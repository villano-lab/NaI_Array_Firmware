--This example file is for demonstration purpose only. Users must not use this keyfile to encrypt their sources. 
--It is strongly recommonded that users create their own key file to use for encrypting their sources. 
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
uWcrLwz0/pgdhMY8COwf3YCegqM0RtMJR8koF41uwZpXeukhYx8zSveMkQ2jfKOmD97opkwyuUa1
PR8tKij3n+psPlzcrDFTiUWmZdL8CBS8vNBd0YCBZbiENmqfmqIN80dwDMLScF2fb8z2x9tr2tTS
6d/PbXb6AQUfLNQh8b5QVkSYO6dJnw7SJBeDRjUIGAU6gOoiKZzDodyRJrPe+KANXGawkMKy1ZKL
i2gL8GyIYkPu5oo0Fotw6oFMRHQ7Za0/uhqxpNMl4f/IOvUMtwhvtSsfJL2I2h9Ow3OHzespIaS1
VPN17PCdadybj+8wOD/RUEW5kFGmS9iVjvuGzQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="WqPbuVWmNs33lmpGcbIxTTOczNOzPRQji04Ki0bFnqg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15312)
`protect data_block
xeMpx4tVPBOa55/k+IX02EMkFHhTg+LVgA+Ftw7yKgoNwEMkTDbVc4BGox1vXNw8oDEAw3RAB9ey
vJq5sZytjcaRtFgGiTKTdhCU77+cFheH0sXKrb8AFpvAYhT7MsppIPuPL79FM7sbcilEsiOGuSYX
Y0n6Eo6E1+QT6NZoXUduXMzqLQBOQmrOXSHPSSAb/lR8rUudkUfkIbwpyYRFPdWg6vKPV5RnK4Pv
pw9CweVzwVUDB7wthZpd5fzarm1ye7A23sFa0lJ0QInzfhdTcefvv3dWDONqfico0/S/MPmxLrJ6
I9O2Rh6b7rF/od0Wxm0rUQI2QXqeNtaMn7QTLVMNf4jkCW5YbSTgnuhJxQZ1MeY4Oiw3m1eQm5ui
8C1lihghPRCndaEfOFORvMTqR8vddgAul1Oez7n4SWw6bVsjI6fiBW8MVYBH5pSHqYc8bPVaqOPX
GF1K4nkspOdYYLRabEks+beNAxAsS4/qS0WrosUjZXXanZnfBbymdJJ9KmwoxuA3PBGpBAyxta3U
sP+OE4lg8FRdf1DvPU8BrWaDfny+9P+pkxRjoiAoYbMX3zyoKtziBthvHV3Wvj4t39HbuGQhldsm
sg54UeegNKpQIzAWx2BfjTOEOnzJ4rhmbMBXkfrqRy+2FLPCK0Un4DrVQVlpdx7xW+npwTULC91F
1KVA3+FScNL+jhOeaz9yUnzSrcZqMkauBWvBOB1fRFfZiOCjBajXnhN9thzwJ8ppvVf4u2DeH3Xo
ew+u1qhZwFPfIsRHRXWJvpjDJn1TL1ynUzb5e+8FXykN513B1/CAoet6OxhSspXrLC4RmIKuNGJ3
IUzq4cKJD1sSv5G6r2ipn30kE2/FkzOG8xP8e+12goqq0lD4omLt0MWSgrptTQu8jRDR93tvHf5a
Zpd6ERyFN1D54zC3Z06j6vFwl947D2viSn/QNEL0BSR+b2CtEDPUrewIllWd9xR3XiXr2zJExQ+g
X5ePpEAJDpJZgzjCuk5g6FPcSoTmzV/A3+zP8avfNF0nyWLQZoVkaQeHWxDHhA3qE0CraZDTKBDE
VZja9uIotxhNRVf2qBfvjW8LWFDCYVDm5QsrDjtQBNwJWYPNsulwQ3lc4qfb8tabmAiF4FExn32u
6W73OGeEHy4xBrGzfm5NRZJUpOfq0rE9QzQhroJM3bAvcMX64yRkcz1FzEvFOE5WN/gEpTWPZUQF
oPVY6khG1sJkHD1BMBV9gl//DwYVx1Yc7C8wT2Y2RSP291ZcgKlz/p/4HyeXW2mUdZD4V+QXymbr
tabtmfGTgHquYAgHKjglRXsLrNGVjXcsalGC1KWycl/XevJOdmwk2nsgdDREKGm491pB9VoX5lQk
lDdNh/4jhh+RzFPakQQZw6SZJ4zV1tY3HggDICPxCJMBGE1KLgOOc/qgBaWmrL8VmE2Tf3UTfXnD
EXmZ0u+9AWNTFQA3lsjRRODKS96fOtFrCna8A45NtZCYmf2j8TOKCFTde58evqn9ILnHtYkwazBV
s0xORxiEje7dwmG8pxWZMz1/2lrCGy8jZ1z1GWN7m2xEIrBRhM8Ts1gjDbj4UL/dK43SNlyRaJAc
TV69IPUk0glsvxvYf9qnvfkFdxrOfLzSlwkGQd7qqEQ4AY/VTiM/6OAjpnw67cQ2Y2LfwmAwpJCg
BBplxeRalAqA7M/1vBI81SVCDSbWkCkPthNe7yfWeq9ynl7QHNWMIb6PjUxnmlFEX5yeyOwvijKk
UT62Kh/T2sdDh0ZbuNNg56zZc+2Aqpc2aB1CYDtSY2rCHPtAqDSDgw/K0dPGLVTgGFTLLssCRcKX
S1KxupOqyi2hvFAlDkNbiAyScAQOPu7be6DsKFXBVQMU5WUI49PfqGyL3SUlnjr7wDuoBR8YZOZY
WcuprFLZwioFCxTXuy31FwU/1YbOrbJtDqxlPB5u9NYViC7Clbcf99eM0XS+obwZnpofhkhtYD6X
2BSo0i+GVGGcglboMJH+/2YyAw4pKQ4xowVJozjPM/YmGK6JVNRzb4N6M7JktfWpEoZsx1dmWRH6
dvaUNmQR7bjmAB0HXnZS281OeI1bxIBqjQgUG5yh05NyNNWsRNnVhVAxehdJj6aqGKHxnfs/ZTD0
oGuoVuDPkG6K/OCloLkaQTaBwzN2UoFRrnMS1Bi97xcZsy7gTaOWY6FOlh7bKnRBEmB9D2Iv3/R8
BzKukTdLKly/E6dxYuAkQE7jOcyyFPkjdurxaO0/akXIC0Du5+RrsrwYo2KapFbb3PNKyV7l9Fly
js6sUhYkDF/TFKoMweVGwiGB67jZiQT1Q8qi2IQOBrJctcNKrv7SDmSG5CBHGrLEjr1Ie0awKbWL
LUYarH5dugJWbFDPy+mGvJyR/oJhTbMJwyCQ29QF5wAwWg0/P25A0nnJyyZoYzhtcZIkOZshZKIQ
Hr10VpbGyLu+YTecASv6SIskCSyNwSNe6myG+AsKi8Iexkc8JDBYZgKZP28Adtjs5tP9yyBlRH1W
IjnycGPU0o2jUEk6zFMPAuuSGurApVMKv1y494JmufLtfH4KWrH1aCQ4hog/BFt7ezJOzuJ8vm9+
cXzzRVa9fCoy2tguY4RizUQqaFRLC2k/vYNAfh6yPaBLefhNJv6mKyOitdQ0KpilseCvRY/UzoA1
ts3A2luS0JLP2vpf6NU7x/Pj6QxAHjKWzHvY2d863A5/SqrB8aqn9ssyjO1xsKu4QNMEqTLSBj4q
9gzIbw9FzbuvvMpgWrBTmVgHb2OkXj0/f6W4/d4lhS6rfiMienX5IPTXwyspUoF96JVGsQMr8ASH
UdO85TmUfbr53BGi5y/Qn68SeykXsIEWEr2NeTqHITtxCIN3XZaxEcSKVLBJM3i4+a7lPuDGwZLX
CTEtoLuR0SORru2vHuktrGve/Q0CIZ5TgndZlBbWGa0oNC+et1bUH3qp3G1hwg8/9mzWFz7AGiRc
aMHo/RWd2qrNa0jKrWX9m+gOBOQDzEOu1AQAScuZ20tP8rykMcQKznQWAyBs6SYr72HcmOumYIH6
obfYn3tg9aU4RtSZZnFYoGMFmXQ86J9IScGhbv2/uoepoYkmr2I47n13ErPp6uWu73XrI3ree1xJ
oIrwRpw33zUHkFmiNgRpSbYW9FTD8jkHn3GPQ+7CPDEvz5v6ZHnxXX3chuuSyNBFmUuSeukJJ8aZ
slPcVAeys+puR7nYeJEZfHseFaOh+zEFp2QAs7rCOsc/qZhJfVRgrJi0gd3GzreG7JKblKhcUloe
It4ZPYffvsypSCSGw1oQYcNqfOivb5ZY6L1qfherxcQ0JLV/1N2ILmD4YlVeska6m0l/tO1YilM6
JZzTg6hMx6i8wdO018B4NOYyC/Rg1M+YlB4UDTJ5Bex/NeZUNfCOOFel8bN3XI7IDutuOm+UDYZq
qm1y+ds7QBX8YstNdZvfrgf/y0eEkYVn0omISAYQq2928tiSH4xeJ7zLrXKM/P8ZqPl85NEPW+Dk
e3IVf1XOhJHLv+1p3OcEvgud31b65jcxusI7jeoU/n7sA5mcUrtc6y2GGEObVyg2emPvFpvfRNI3
ylDPbdjxEclXYU8j+yy26vkN98HP1b5m8R6Kmy6Dn/TZHlbwEcKB+5tmqEqbalME9i0N700DxOkp
VGxSsH4kUMsLapy54P6+l0gbebnXpS7O1DFyEdBUSLFG2zET3uVBAukZocYdRyx7fObDrLfco6a1
r730GG6gSI6Y40LbG4F89xQjQGDAiP0cktElyeT+szPU1R+xhVAtCIj7m4KO2yP6RWuoZBlIXQ/5
6H8a4OsYvbt6hzgh0XjMxmbm+FHxirab85MwdjXnJ5iA4myI9cMRXISEY58Vm7JY5/9Drv8OPzl2
3mkG9T4js+GTd0G7zuvK0/XGcGCyNApugoROvEqgvO5Ng5pv34VMmrdUEHj9VR1E7RBvHgN5FaNx
uh6AFolTrxNR6YIr4EBZJeseppGr627vFn80vkTZQVXTqej5QTLx7JGj9pxVd5YTV78DN68rdTUx
ZT7BLaBCRcUTu1R9PYeVq0LQKmoQ028hbzgcZOGmplEN0JZBfgDNe0rNRvbdzwSoimJJAipz+Qdt
y+zs/fZXSQsRdqXXXR9qjaSwJ09tE1+UdFlSHmDz9jBUxgI32+TDiFY4nABGQjePqruPLvrBs77k
EUAr6MR/y3Xowetxh8ICfgQiMhQuqK/dJfzmf30oupw9ugOn2ZVmxes4AoMwlUhfB2TsHuDjJTJb
EJ0kV+oEJaLZQaEupMhLM/IIExZ9BFMsQOsr9tzNHEftRUys4zf0uev43YgxKn+Ds/FZHnyY6n1f
6GpoEtbyjyBhJToPod7VchdP/bJNzVkHiX0+s52PWCemcVTedsDIlZ/Wqk7w5VNuw6s6OCq98B91
VMssCX/iDyJ3sjkqkX0Q1crxRRB3MLuhxD5u1F6uC/XXRzdqMqNp+oK1AQkThgcI/BNRH4vmtMef
j1A8B9FZb2MNGXbaVcHQcjtINpKTQ3EZ/wCuUZWXYvrCKlYyKD6EoA1k7DnzR+iSA0th8kDuMLC7
eIffrdwlHCYL/MaGkG/srUSYCubhtUs2WO07F2lPzClWtUfiqS1SuBcP3uqZrKmAk2aXY5ucMxbE
tCRtMXRe4pjfn45v3DDUB1vvfvFpupeeSZMB+5gF1gk5JCT6LmLhh2LqbaIoEkip6/QZrc87ITK8
5CsmvQyafwLY+hY1/4t+eMG6Re4MxK1VCxZrtLTP2gpaGG8EE5WCx1LQTByY9qVyWWxj113Z6VRP
N3F8xUMnyGKmLGaNqFiUMNJ+5nFXwHk9n9LEkStpxgfIGvrkj0eZ4Ys4P2QRaOhDN/zjvckLtHhE
eAqXJ99S78HMZuFYPa1UXt+ayKKQqlHdlQF5IRVUbgGrp4+xkW3ihj5JbtzS+P2/LmlPQN5pPXcp
fw/9wDx3QS4CIauQb2SsPkaTEe7iM9ks1WA4yXEHOx3LAms0vhqxPXElIm0fqJf/mZuO1Wv5s4zH
kiBJBtDhEG3K2pMMkYFZAsKyc3AJHeEW+0ragtN7/OyqP8fOYFMWDU/GPPcuuO+CRyMCwMmE69Ls
zhXGrCqHErZaSzbQkFp1+/uFrrOs6kPDIVNHorDLw4Kcaa0Givr0F4Jaw2EBIAlI0X1e0AyoiQ2n
Rp1gAaLTQvwqIyZkwNZAA3haGx8Vx2F6RPj1OHe65fvdqdgUwVzhe8iWNUox4ds6+eo6F0i4BEUh
9hvp9RbIaeDfrYBSjpoK04yQSFlr+vyZ1JFTnshZgTInuVv080I3SgmBzgtQ3c7A7BzkaHgj+OEF
ze4RoJGbHwbIDkWkpRO2820JfASfPekJHF+din5vn3n06aVfz6SrDkDaIAnKeDm8CsYuYa+ZI86I
9EGRmurmRFXHwkg/O2813a5LLsG+1qf43pNMLIMvBNhjbuiPZluenpNmobHyU094w8ApvR3EwYdg
98xyKpmNKtY8JT/LeG3ll62nohRsQELbVHvECxojVCtMguWXAPiXv4XoBpTs/52TZlUJV+/BF2eD
uL12Hic4A+Igd9LWrblfhDqWfTeB4SbuGd8ZPeKDy6VZ3GJk+chQNso341JkqqjFOvAfxY+AcZsE
boBYqtlAENn4EOWsRfgHja0XyvDLKFdK6qWfRTTNlbqoAWD70E/GSd42xcfZnJOQl2CKaepBeCv1
nSAaX5Fp8XzW+q0TCkix4YK9zUTO9ntc3/Rz6vmbneH/8TXI4eGCUbn/EzUSmVXCt0Wqx8kMBpYA
k+ti017uX9z4fJZuZAww2VlWOPdOcn1O7pL5Cy0r5I7ELRkZgrE3FstgygXK5XKhe/CsDdhVsOnE
LoZcgFTuV0PKazlpYedhOMmThg11kTJebQdyXAUPcDb3bTLojy6+ImomHLtPQCSnLtCNsBw/w8RF
TB/YpLFGHRhmPRzuncHYfJfy6+2l2mT/03U/tXx6O5ia/6xPvlnY8d1YSE8aBHAjr9GYHbuz2w4G
3goo69PNkW3eqFxzgBgsaAv7Iy2OhjVWU2zfpeEtWqaPPf8G6WWe2vvvbDSlMyTWirlqShQ1HJjR
gyBE7S5WvVZHcLeiDLb/LFyDjeCVQRrmUYqeIubnLmQfqVVs52ESzFNzAPhQygNejGRmgOtGJx29
b13q+AIS5fRc+Rt8kMlGPfDBcqu4pKTDB/M4uevvz4tsPY/rzCHtqG/zbOZjo8XmiyS057wfyw+6
NUNAcRRsterxtQ0E5ZpG63CWfK4JcO9nb2c6MlQGLx+kpOho703Qk/rKLBa5o2tQl5EYExH4pcCY
Vwc5NEmLx+m2l/wZwOHJdEPqxUwMKuqVcPu+rPJWWQ2viavNuI00G5qsIB0NvOzwxuM0OAVEK/6s
0U+bJetGe+nnUVLdSZSIE9Y6MUpLlVJVB+K7jOkKfHfJOnN4BpPNMhAZrmG+hXxNJWrzOzCfnrfY
y128dmWcGWcm8sfOx9T401rkG6QCaKvepQmGS8YXVASBe/9APrSCdKu+vpR8l7XR6/tSdcafVai/
pU7wjWPx/lvsyHhqoK6vMm79bqolGagmBCqEUVo2cQsmgfA6DcdG9R6gOIZRaO5TpsWi809TD/W6
w7WF3LN6W4Fa63XDuGV8OwrIM/9QeUB6zQ9Z63wskTnJ8479TJnjB2//T4rTxfmFPnkRXI3Ziiy6
dFo/ftordh19O9he+UQ06cxUZSwBXHr75GEjnCJAo9wWg5sVMxSqcvqNyEdzsc7jo/oai67IMPV6
yynmQVtr/OkGT4J2KmU3MRj4nWHX9YDLkaqDUTqKqmWMKXDDZKAilHSLZWAAxULSRDQ+zS8J4GHR
wbMClk8DOXERHTTyNFQwDztnQBm4OHffV9orUrNZ6EKWNaCWC+LHRVDOSZtynPiPGKjNNaKm9tEe
UfNxTslLRMrnl+0s2/GSHZJ0MXh/ffeJp/CPuGgSYCMAP4D0nyWdvjqIc6wCcWva7rzDQ5aBjr7L
ixu/gVT9RDFYiFUIM5PDSdk5mj3KBRFtMo8uAyi39fPckn+75uGeloVES39HQZUsP/bUHwRwanr6
yQ2bhn+kRV2t8mOAYWguX9bYbIISWiWQKPBvHGVxF70FJVijz7Ti4G3Ny1+ppxE6UA5nF1c7r87X
ouHE8dAXKpAi0UlycyFY97lIHX9sL6Bf97PRa7vuH5RIFOVmIULtlRsEDP52or9OEjpeEYOGGtCg
mcQy+HyEenjxs1lnvjMdiumj707EWUX8dfW7dkPMLA9xSzp8kCT2b45tl8IZ5x+HPrC35W0NPgFx
+z9fYqLZHaKGoYp2NLRkZdp8SDBEFCC3vCR1AXeqaeqH4SenMqElanb2xQmll34Gpx6HvjSPX5dS
+MbejT6niPrIMStUCTU/0CrAAG6TvyxA4yVncauz62BpZ6ZNenSnh2dWWaXiftqDurXkUwoBBL6G
1QpOAulFN+9eN65enVSSGjMV/bVAofL+I+bcP0NCcSjkueihqasDK4Ro7hpzEelS/XnVs+I89Gnl
UAVYoSSTudp7WWTfFZ3oOppJgKtjtLaxpM3vNVOgZmE1EtVgvEp4OR4yBvs940IeK+sy9bLEnjwD
GAkTygz6GnKhK3ZFBNJvXFkoVhoHEJ6HYhIqKWkFeXekbRC2oTc7JNnRfB3D+a6fSP2sTdyLeLHM
qlyDpNFhWMgIDplmU62KYs+vePWeWQ9blYaR8GtCJRqJl/Ka1DehyWijD3mf4dV0G+eWP//OLhkW
DaQwbO/P0+vVOGO4wbWr7Q7A83BRUbSK1+D/A9G8yow7fiu+lmJY85mR1sJgaz8jyx6/e3qzIY8Z
zmI4boN0xwqstuptxqcB8zIP9VkVUr1VxAClefierQpH+BPVby8+PneofyOsXtmTnZ5omkWxP/fi
QkIySvn0FV/z1z/eEjelyW+JuHkmZevY6lLOavcCdCebhDDMCwjqFxf08wDOFqxV/RHBLKkrMVsL
63A1ET0fHP82tfu5ITs+kerX6PFa2px0yvvoWkhuYpGTImeK3lCOZwuPQyT9hxFYalRVGmUM/N3P
guk8QH2r58rBaIhfouNugQXrz6HXtAa4KzICygfw5ADnruP9f/rr02+xPG2Xd8ttxWdoB2l4WFOo
HUTTW3EU8FPAlbD7Ul3aZU0Rxc9A4XZbTTmS8/5emyu1EaWtNaJTL3B6zNAXWpp3V5bKArAgs4qW
0/wuqStprLiayhPIHGgQOiCqKLRbpgGCNQEXgnpFic9gAdgFpQVjOgFcQlWXTA30whTc4ylTtOTE
sW8yLw6DEhN+Jo190Zeyc5JFRqOX9wobbWn7FTQttLuWAHHHBPmbrcw70r9FiVim9ay/2Efo720C
E3ZX9l2JbFWybZX3a6jME50YJb+FI0j3vSaI8PV3TEdOAa93B674T1eY90/OmxbtK9oNapnTmpgs
f2DOKZIBM8v8k9hNk3TTpJ/jgKJzWlU6KminUfxUMJWsfIK3eY//yDigH5g/sPrhx55NNWP7ZMAQ
/ZZ9DjZAoPHigkBKTonagdEXsDeuUWv0X87hrCtaI5X9APtjcSyDpDoaatnXsUPc6rUB196QP1Oi
3N9RVq3LjVktJfJxE8W5ftFm6YG39Fp//425cS/sQV1VHNAWyV9GXgjs5bFmPGHY3BHCC6flvDs5
y33PxODrMO1HR74PIxkejM9/bEGcwNZvRZvEWsA2xEMbidArOqm8yobYzJ+LdXV7RjvNt3RSIEHx
CZAZ2WBv/cCxlohByEL2T1e08jzjCeMpWt5FdJJlhR+hOV8tr+SMDoS+UCRgMVUvobkZ5OUwfpxw
vR8XMk0ILZFW49LJ8a2djB7tVxZ8hiU1u8Zm1QiyocEBulLiWGLGzY8vdoa9wVzLfmmw2W7gNBNi
Nc9YGZCCyU2mpwkCON3fgp0ohccdya00Np5sB71W6ANxLt1J4zfMNXvZfsH97VLV9+Vd5NpyKMgm
SdNUkggv771vinG+wk064trAVkmIEkQ+hJPNJkehVz9vxvee5nWaZJRDnRgDqmTxff6nS5e5gJYU
mcHuTfX2IVClXCdmVzPRJeDOMdfnm+NZZen54eVH91zEWMFjN8fJ/45XA4oqvxbe3o60f7HZ9U/M
5ciHStHLylXdaRks+cVaSyKa87l4DPgp7vcZsnEgvnvhGrKOp07r5BJn1WCwBvVn5QlqjW2w9luS
SAEnYI6LzkZzJ5ZrOPgX9wVfYudjN39NMN/C5iVxewysma/j3DPvgYLOTyDTi/IDw/GqFh0MXxCW
xgQ1WMh3JlCcPA0CqyLtQ0uzePm+K7Ek7krJEA+9ixPG8snZbwoarhRoGdk3zhOX04XB3xbG2pP3
rD+MzobcyvJlVeHhA+xQMJ2F5EoB0yzCToCcq1KLo1yaNMHiv9ZfVhjetv36RFIffHUOHVrwh2EO
uxRNVOltEMS1hUEs+Unxpjndi36qvleMoGKG5SjkUWrPdg55SUf483APiEKrDfadAtbB23PtU4R6
F7bcW8K4vq/810FaOVBnUPzGKN/tDGtPP0q1FmwtWDJhh1Ik6U+C8uDcVPI48DS5qZTOxff4S8U7
22lnu/VuIxJOQ/WTaBjMJ0m9wByDKvDxP/ys7kS9PdQ4KT7k1MpBFrjDFn39K+7B2ZGLNv977aEI
AdGtWWeairVgGikXS/CmZbo/My7IHYGftTx6lWdNdQ9pNc43bAVgV1hhQHmp4TtlUKVD807hw8Tp
H1P+lJIZOW3xZq4Z1zZlE3ew5kzKbsxDkK8T/B21gAqOSZ9dM9815ttmL41MXB4U5eTFwUvXAmwX
vPSotsa1XaKcxiPalbgdPBKeHbwunQPvFfv8TradZlFu0wJLwIfDlmFfzLTdNQQhFp/q1Ch0ScW3
x0aHGLJMZUgixA/RauOfTACI4AUFEpYlxeDjH6ECbQ7no0B2k4xHQmLwFB4nom3s8xvAkCtonENt
rnf7YVGLFkSVU2fjl0i7yo74kQrg9hh+8tI7FzZd6POcRgBYq+iSuFgnEW0XZ06gzB7ATtYIAxU9
7n/npJk6zmr3yyIFH8i426d7mxxsVZ1vGpT4z/9CvqDsCwGrpkULaKZOTDINM600Vg6oSLXx0a5Q
usbmsAZaK+ST4X+P/B5n81j1UFxiBP4CGbYn3Abbk4S1NHJ0TExJ0ItqScdks3bcwPk0XIziCLbL
t3BmwBvrk2RgH6ZAvTSa779R2REvMpyQ+epph6fIFGauobv19eF5MjaWXUoAyQpJIgClVak7g+oI
embzX+UM7w/3WO0P3A2gDpme2BMpQPtRaFjS88wnEA8VL0vNRrCe/oRKnX+ZcxJmbQavFXrTFnAV
tFLpIjMWX14RTKG05NouFRFziZ+7NhA1B4sKHMvX4ml2LyedMDXVT4QYjBnm72BNNR3IdKCrY1/q
KAWlpDUwieOGD1tCYhi//WSqq3729uksyuFQv+PkhIIdqAMVsW4nKA4rRWKf8LF+ITNZk3PXBTsT
mweR+ZQIx2UyQaccBmDrOkfitTbkFqiQqPqYAehgFN3NmYD17208eWC01Pq48QJr2gazca8l/Hlh
3Z4xin1/FpX41e5ChDQK84b2y6yi+8xhl8IaunkZWGI8hXXb9PNf7k1vpYN+HdjhaBXaiNEu9XUM
V0ZFQBF5874MDvSL1GMDr6aaLhR9Bpatsr2lCH2oTNDn6e3NwsTVyiUAdD/nXXMEH2/IDItXV+ir
vcCsvtv2Brb+EO+fy5S+Wqxifi2xkp5n7tp/Emqkolq/EyrGAqy8/q0vu/ZydkclmXESg0Oulv6l
VHrSR2WTLAkaIgwJ/3GBHQIdI5b2CyK4KzRI3vUL+IDicgWZbuEROplQTFv3GysV3TaQesY4iIF2
LGDLdfk4kTKeiv6bM7YNZySLvS3n4O0VhsXgSfX4L4Y2TXrnAPkPzzayLbRlgJHCEIdCsJgrjlSD
d1x4X+ByCTvv1wWy1nf4VSz4F6SF0JFhs+ZTf3U947RUkT3GIh5hyWvYnz/B0i+F5bbCGXjy5YcQ
W8t5y25/4p98TmWt799UdIAVD+frK6bPV4naAPKDymbUBIU+/rNup+uoRrPnhVSzoJKAULCg87La
o4CEAiiW/inTA6kCPOwQqB6DUlaQehxyMbCl/9lrhTQ8BqJfBuiLW8nHJz131zDibwDhSyFNBp2p
VUzFHjt/7mdLXasC5arYU+tfds8+oNP1kDhdksjPirYKFyUKTBckj2ZEqIIJtOcw5ISgGy2aLBFY
ZseUeXiyF7EWD1UMplAw/Xf/tU7sQRF2U2qMrfFYlW3pXpRjlIZWzJu8OzWL5st49S7MoXg4Qx71
DkyCszABD35wnfEHd5KYmHr+LrSzh6l+5/4RDLBIjHOcBbHTBO2MOasKPL4dsC9uYxeqgakhiOW4
33UfppQLOIIjRWA26XOH/f+RCSiFpDWwoHgiRsSA8jvvNGrDeUaVhV8EmF3LBAIPJiHZx7/1qUlR
uMVZC/PDLGrfHyqGz0gYBXzisXFn4JWeVF3Q6tehdT3RFeB0aTr2xP+I+5Vp1iRbaUYsez9JUNnz
QcFGyeYVH2GMEyMdSaoPgBEZdUEf6EG+Mq/ZwY+6/DXRz0JqxjGDy+X3WcQXOcPEK7U8qLfp7UgW
zgLKshP2LxdxMwY9S3ARfGer/ns0tObCK3y9T9vgPdZKrG0HXYQO7HI6M4x72/3BcRr7GXWW5sdY
70hfVmiurPivC3XppIIh6CqTAPTGaJCgdpc/TzP/x6FLWjWvFUr2Oa+IGN+kAsa7NgsJObuollr0
ypo1UfdIrwJhuQ5heJQLMS5Cj3hsgEWtA6MdDkSJWwvjaF0/y1n5vbwSf8Vgt/2m5F81pc3bbON3
HerqGggcEHpYEDQvUDlNh2/E9jKKhKdWDORv7HKqtUqYgznIhoiMq7HCVc3smhXzi/JLNXYycIhl
PhSEQhYEVL9f6UPNhywdLR4Wb0P2WXLrP269/CzwJ+W6fsGn+gtLo4eRQPCcolwPNXHDzL5Mp7Bb
l10CNf22HDhnSQ7Slcv8PP4OOz8GpalCUPSxyjJhXF+b6vxgHcDnf4lnZHQJVBlj4yga0DlZZRCH
OcBr5f+Pb+//bsvG0lijqHIaCuPbLqqFi5nUBHJaqAoBag8xtVxo/6dWBJ6VNagDq8rDs/uCucoI
sndDw9E9zAoSlm6g5ZMu3DWGeVd9Cbe4LJxKgR0uDYEy7jlqOHQfPOShOKEkf1escOqzxuRL9Kuf
/HKtwVI3NBX7sWigSq7srgInkP2NBvAgw+W9fRZG4ANLbWafuGSkeVMsqeEqocoqrOUoBShsj5/P
o+ZAzSS9Kg8F80xoLveLm4B/Vzg6ROrGJWbV3qTgr3u2iw23ZZhadmzDElBQK06kV5VIljANaX8z
BZEJ75RyqI5Yv8CBHR7wsm+6QQteHhjSncYegWarRA000B0EDjTJ5e1q0lvYt/71Gs0N+3nRoVW2
YYlamwxLN5y/5rWCK4tJOFxfEs2uaI4XLgK/dU55tfuZRr338YWHsn8hi0U4Ypd1Yn3w+E2B9JuZ
Sp5TnHlCvuCq7AS0nQeMQtIk6Y9+YK7Vc09MRC8xb3njSJBgXjscvPbY3H28LhOxYHdalCYe8IS5
6hzXkH5fSuh8CVZhA35g8nYRRSAj2cy8cmFOIuGmQUcbYE2mdtu3oHnIkml5NGCupDUCB4qVNm8X
gP6ms97HEmogo98XA2nexoeH2FfRypuPzB3sT1SJmD+dlcQZusn+1KYM21UV7qoVGfM4VAooLnA0
x17eVFtTw6v5gLfxi9fdBB19WHwc6jj3IUjydgajB9JS1QzikN53IMwoHYJsiRUY9UMy0ARPtglq
/jiRTVtag+oy5Yq3RgrXlJZd6u7d6B74vCcqHFVtmPr114IkMVPes1yfU8LTvETt0N6NEoxKHbZu
h+sWyLsn1kUpD+Y0gtzxlunpWMm4nfMnxOIjmtkAWQybd/RyziOEQ/IA6o1r5ACVgMWipwPe1b7l
6Dm6htY63m3KBUZRIHizVZAabuy3VEnkI4YXY8KbjzMVxpeH04frpCUsB4YwBqIb9RXvAP+GozsF
3uHbJWf5mpcRdGy8/sT1K3NL1d9JqkAMeSwPPv5aJKRFpPwHDcsQ+RlSwuYx1lWLhXOlEVKiCDrL
pumAQGUr6nAg2FyK7Iwm1nUzPM+i8KHJz1Yr/u1Cp2NgCKVay3v0Bc+DKSlExlHM53NxhGamDFec
cDuQa9c+uyRNlCoTgtLxNEoFnivm2uy1hzZ+mD1kThvPlHxpqoyVMRNNw34cnSTKHsN2LrdfeZ28
mE6K2zCSQ3UwXFS7FqRbn4bGbiLJLuJyoMRsnJ9KDcAX6KxqbXjyGWCJtf9K8H40NyqnEfCu9CUm
JoyqFVnmA/+rzVYwne2ZLhxaov8HsK/w+XO4jbuxmoTAr9noAq1aONu0z+2KuOLkwX2JMepes7A9
od2qyjhZDjydA4luKULbEdl/1SJP0eYloVFjzPklRieNWrRnHgYmcW/12nTBqf8yYJC5N7pS5NqF
8TtV8sTrh51uFycMMbsvmxciZO0yAkrVEVo4szPdF3FaqdiEUm7FcN0i2qSQzkaQfyhjTI2MP4lN
3rxRXnHfLMymtW7eovbO2+/VkSXXFnWXWSN3H6KP9LkAVFcdw1js/eSCtwevIJWWDNWfGqGWmNgf
07Vm6sJPzHvB4PKEPjPPAQP3Nrz4Mcis2p/f89MZH/zRRRPnz0CstYb9X/g+k9RFThvsCc/7Ubm+
OUrENux4QHTLe03m8R68k/xGZQ6r5u/0OlGOEI+8wf6LP7K/RacWUDp1iqbyJSIgiVaaL5iMkeKH
HDwHQrEcPvL3szqGI9AH2eHsia+hku6xqA13RZznnBSNAV/QxU/aLZ5AGR1Oi+dB4flsU5Ha35Dx
Ylbcn8sDdrR3IGrBkaMFjVV+TYkWLVOrnlfDSAZOS1ZKXofPCYBDyuYE2Uqu/m2dZ0JURD0WTOUy
zjxRYaYI68q+XTXbyxtzDw81ujwYYjvUiZDcaj3YVLUqSJdbaJ8JtmUnF8l/YX2kJAbqcrI9+H0d
f6CBK2kpKA/4+mFEDNa0cMoPdoKKDG9AQn6gn6JH/XLzrvYghXUEyTUBTqEaCL2eQM+tKLa5+FhF
+zBZlv2XoWUTk5MHHdLcjXpX5Pqpz3bLk1ymBLN3JoCtVR/Q3BQ7MWMeF9WbHoz6/aTa+fZ62em2
1Ahxgu7By7NALKBiv+qz6mZgmOzn4G3sKhYNMIQn13tCWMqhFlkMClanGedzigsNAHs3cVSBgekF
gozDqsCVrfVKH04u9IhjHkrfc6cPUBL9pMmNRPe5qRWQIRX/bUGw2O8ilyt8JX3Gabr1to6X2RhC
T9UC8Yo7OwZfJnod3T4FvGaGhAi/wnx8MNjeo/o3y/G/dXQmOl4VMEbmwSZlGBsq4+j+VI2Yw6Bg
H51IVhr6xofk02RyevvFa8jSAEWrxHPQP5YNm/NxsPg8LPXO5wTbJjMEDnTuC7s93cyZ680ROS5H
pdtuFOyoz1i9Uhink9cWT3vKuIrOMtslZCQaK3EtXd0U92K7HxYpOiwPqaw4ci7rIPbbg0LupC66
3qbIkvuZkmSqJNGzRw8L1nNQFLwK3CkVyEI7TrwPVTvitQeCyjchp5OC7gTntJiy5iJJkVTKNJJA
ZlJe37iBP6jVT/rWIiWdaFk07W2Y5U5Jp6kOyRQ75sn8erQ4S/dtSklqtmfED5V84iwTstk5qE9e
5diob0U7QYh10y4EHaLOqQf+ZyBXYkm6jdMYDhYKD7hJm0xu0qfjIzR7uWc0pESVvTKBddXTCPuf
HMMfnCMzeKKIHwltC8DP2WLfLiRoxXt0dwQypwMkFQtQSmm1/zL89Sc55yPlPgYvrYv3nfZ9xJsM
O+0VgY4gsU0nV/2OQJNawxt2KuV8xT2xlZnLw2QlFShHyqU9LWo80n8C9g0K+qP9U6ka3jmxl6Vs
n1aFOFeEYF2+Nphs82xlrMlpa5sfflY7S3Wsyl5tK0Cu8iYDgjm0PXonaOpmYBdKJj259D2QqUet
Wv+afRQHO0tEKPgn3l8ifkmPznYQhzoV7XwB7oqOn1lTFQ3wXhTDATF8itoOFRB6UuI6JlEVR5og
nOKnrVLE95COooLyt5HFTWRUys2oRd6Oh/L3WIK61YZHpshNRjiH38dNbCAQv9RQ12CZorgEo/P/
sRddmwR9J0LZkAd7rit6ySArmwqX2QmkAFCfnHICdTT+Jr966xVAk2U4sSIqB/TGqj4n6CVbEmf9
3L30Zjv1CE5ka5klAHYAi9ZjBlXev1hCY6nMA9Gxexg5S295ADRDU923fbu1wG+mw8vd6XdWGfgD
WVfFaxeCp02+IgwFX8cPd8iIWYrJAAZmqGZ4+CTuEqvnGQoyBX0clL5F6NEAmE1Jdy0Z86j+Ye0M
JKnc05qfHhQDLOi4TsXQIoswAe5vLJUY65N04GpSSgIUzIKvS2c7kPDnJxvhcQIIXFEnl+CBvnDA
+j2eYFgiy6ZKAHlWDgE6E/6pGjHYumwSSCtesQxMTd1Ale53rDvu638/CsaHxqv50SQsg3Cs0r5Y
Mu+COYVW+DH0RO0p2yAJYBGqz5a8HEHk+5ATmhF/0ifJoNlByeOpZMnIfI/XRqy1zy+t9wY/NoTs
GMI72IbhKTl8we4q6HK/yByPc0KQR/q2VxK5qbv+J1s+avWEsAgSo+ec8Ehfh4prXC4ByrjLG1B6
1H0aL/2AZjhcUwWdV/MLxg+QtbCoAjD74H25SB55hCR7DVJmXNMKhJETIQw78aK0njvQpRmFLVon
UjcyfW+tdT6s5/H9Qwt1lWJx5W+Tc0KNBSmD+oihqok1dBSf6rF6CZ/B1EcywPVdNwVnLzJXn3vT
J2oVfH6vV/LpLUAUy99XD8xS49e2eVp5NiRgmNhKcJvLT2s88CXopFkvHVj1/57lGmTbqnfOfa/F
qMrU9PLqqZo/7TyMhso/RgI3sSpXMulBceyamvgHaQy7euoWJjBeF5nR1/xPOr773RViIz30QLAx
U8EZ80dQBu0N1pm5cikAXYti1HqaNUpVNTepjw/T8wm0LZQG7CPShYJzm+sMjHcyBpgK5OhFCd8T
/GBqrO2PY1xaVogbdYDH11W+DeuRVU/4a8kOndjao32g4n4pqquLd1dJSDZmThBefqUpg9mpI/5W
ZHYqcS2JNGT8TO5TknIUgG0ssib8bZA1/kXLroaVlddylr1EncXSV9RGkow8ckLP/FmRYZyxc4QC
CvgZFGhFQNDsFmEtFy7NMpTznu0wKx4ntfP+OoofU4W/HTmYVN/h0zC3enqj/58VdBGWntZ8tIF0
m1mJy6xjwp4LDlxodm1skG2XJGaVpvJbfrxYmNUUop8n7eBZVl/GPjJM/2dp86txkjroa0bHVCjR
vJMFsKjg6atCyp3VmCfizeRJEztpPvChHPRfh/o2BOgMWXbofdXmeK4+IPCbigP3lUZDYjByYQWe
y1OckW+6I63UG1+O95MVsBFZctQ9VBY3uBHF6s2SLanrtJKcrDf0D5m8ahJcYCFT/5lFe95amcQy
uf1Hs6Ssk7yd3vi7FsrtNi2r06t2e9o5w+JcRpmOV+V3+OPPiLU1LsApcCqXoew29Jlr2R2MncfP
IBwDVxS80KgIMVg9FxUzJ07qH58envUD5QbWAgARxEDuPVFHXumHdXrD0BZCenEH0yTiDe2RkbOC
P9qDWEjOcHm7RXa1JTYefXZ66MVWAhBIai4y+342kYncdQDl9w8FT714GXfppbmmC/RmsFWFpcMl
V8ItSQiX/Se0nhn+lY5XfOAg3QJA+WAyWshDAV+UAt4V8/zZxc33+EXx05gKSl7CvLlmU1Vycno0
pBs/Ih2MOHBEkPY1wMTPrJSFgIejpbCx7ZBchXB9s8At/N3AZCMGmJ9BIFuuukkBHkn04gsP/pyl
YZaKd+3rXmy+Vad/p1pPMFczrWCXpjYHklX4qctHJaAxXx6LFsOr+wgWbNcM11UrJhjoq+RoRJE9
gTqCIgP00/wYtIgIW8EhzLXac2rTDm3ZpjVvv5+kquBGiZ2FC6P6nIGZ/DUm6ZGFmCDKansDjCJJ
1TDdHBAvcV/NKnpeElhgk3Ged64Vjga4uUjZ+3KmKAORfVRJ6ULw0Gb7A24jYlNBv0oWguodUCkv
KuqXw/G9y01WJ8AsWnccvf8ovKnCOTRt0vDTKyhkCT8REMRbaxFXhxJ+8RNWizKWxxG8dbR0fk+F
oYommp88ZGz5zaSAB+HqWOBXPHIT/fezGyI7wtUoLBvr1TEYkH0Z96YAEp7916amkwzBtibJ63Ck
6VjgusVy/7sFTBGo4Oic5MNYI8UBEpc3QcnrtQKI0uVBxg2ZZ5Vm9jIAe1oVu9dbgoR7i0/UGmyo
HuC64u2patjG41S4xuIxZsu+am7YGlssThiFm8R0nsskxnwwUI1y6in4+R0/MgjD16O+oPYaveK0
goW3du9qE7jXw9TzCykLDqwaNnStailgAr/a9dJ54NpIXtL6NyylYugIf1VqV6jNAgFM6jQYhfZT
5AEwMLus1GWc9zrJQbnE4C8elMhckp0IOybCj/zegyPNR27gz8tD4aaa7YiHvG3/ycPReZhVe/a9
aDzDp/xjGguDmOJlmTna0+HsLvvpoJPwCUqoHrZLcQyw0U/whkk+ph0fUNCLNZKFoxn7s96SLlaB
yT9PwXtTYCR38jv8y2gnnKUwTMM/LivRukYryL37D64h7og1/mLdYinLzfr8kHzL9a8dw9qMsAxr
LzBsXMJdcYKSKsMxzEyO70DXvXyk/YU+SmiGiodrfWDMbaIVjkXMVe3IVCmF74RCp85b0B/bYn6R
am71Ix+l8VKev+axHdxjuwSLNLNkSisEXZ/5D31x0e6U4IM8rS3fDAZ7GEAy1b4822ynQSFnlUqH
9AskYyTnv0EsqnjqYvy/EBnnInfOcSKt6R82UzeMrYn3zoxLU3zEJuoky8vcaSmC1chh2Y/YzLqA
2MhBxrQSukv5Ecx8mXFqnb9TB2ovPToeT9ulgOpk3r0P1vJ6F0mZ0560EM2EPo+J4OFdoiNqtNGn
U2y7xQJjfnBkJKAuYSxEgjyJBFE1yJu1i2Hmb0VQOW+uOuLCjwRxtRZH5VkzIVZfbmstGLrk0DU2
xaeGZkO+ZcAhTNO9lemqURd7gWm40CQsrOo9bodM43WwI/fQc5/+bmSmKYPiyxwYhX5TbnZzTY6b
s/o8F/Rpumj+j8Q3zyHaPWTL+2vbnWkcml9SSD7mWglx5qpKwBm/6dFTrHL3H9hc+YRChOAVapu8
CsobDV6hbdrZunWq2dwQ7nOFJz5v4M+bJyItde9cgWoJuX1VdIptO3tRDPoASq6KEsU9whX5Q/HY
gdrSvgP3Ur6Gw/5OHqZXmESrw0+gt+MqEHvK5+aJCbTSwvFuvtO9P7M4BB8Hc8/imh/OPDhhnqq4
fpCTb0PxsDQso+ATAPgS5zOZ5lQ5h7kgNDRldR3pp7V3bT7gFkHwEuqb+cWhEPSI6MrqYQIbxRJL
Fshebc0NghbVOzGo1IHwUroxLVMu/0XAOxLeirT70jouwXudso/+FC00t74RahUKR9T+uH3XWmnD
lWDs5guvqv9aCZpL59IfztB90x8fh5PYiMV4+sgtMNNJmixh2pCCr9JAubJCpFRelxnYhCx0Md9S
VaWEfAW7Xrw9NICkjF1DtUA/CNrY1VSVbsA01jFLNRdxt+79YGEyrvh4s7d8sgkoEz++wxS064SB
LthB6iD3xa5C7yHFJmdzaA/4xEau6dba5YG4X1J+BqcGcjxRp+mOlMLfww8pttDi3fvaVV+ixaj+
kjC4KDqxU/Z9wm6Ojn15joarEJq4djYRpcTOu6XCZ1See7+QHiCcxDUTfuboRfBQOzWGRyLxOnMn
b60vxTqgNP5haNhK45ya14iiCrhRCBaM1HpVo0OYq8y8+HWyuskdzjNcUqQYmH7ADaSPEDa3x/RB
d/1O1nI/EnEgI46iE+emc1tQQ5JGBBNr2zZjUrSTy3c3v6pFnUPkhvlpLOJh+/9y0nqDtlv/5Ec7
ZefDiuqDfRTXr0Q9ERZO0b6YNUi1XshRzvjCiTXVBmfuo+NqknTQHtxX/IHz3LJVwt+q5ov266Qf
F43MpIACO2jnhJl1NK0kBBPwZDFMn31C6AoeXHB+v7FxavTzB/JzNO2d5pACMAlMrEKPVS4kX8Hz
mrBwV9BgALtjK/rTRCWGj4tJFKuHlXQkZdk5tp7GyfDcNXuSpXNGcQN48XPzDrM5irl77m91cKzS
09iRfW6q221IkuXfZwcoQxAXcPEsTf/dzDP8fBSJcLrnwS/wUbk2g2vBf7y2xrMkX5rOp2o/KhW7
4SNOCTQWO8ZP6ImffrzOkGrBREcpwdBMiNW5SX8Jpga0vbqM6GOWLGJ0pp/c8zCFwOdVFN2ZHyKd
GFu6ofPE6IH+0mVoFobxy1qNZE/NCC3jmK1O3I9cCymO+fqK3jGzIUvmDZKzDLyMozcYok0wR0x/
r4jBHXY64OCaWt5FKjCXIAS5fBon/tY2KOe/W/UyvdIPFJKgFfHIo+EP7zddGLzep9FkRYbltKEQ
LLRK6e1/GWMolyMQ4ud0uQfKrqVBZUOjdhE/mYE92XdhrjjqQHyf1wokfVQK+QcDmZmOYOF761D2
LYO++M1D4Utn2KiikX7CAUrF0nOP4AIl1wvLw7C8CXvT/O+NewgKOXTMgkRMsV7zItEs5OoIcjda
IC6phjnG3C/f3HjLiIBTyxBc3OJTQTKGbY1aZFwujm7eHnNe5OljN3xvPPXeFKAuzKhx0NV7R7Lw
gJbC3gjFSH+2Y5bqRs5Nju7J7XOaDDR8b2189n/3Q8uTmVy5MHWE6+QaWUzq6QR0hZYLeNX6s5j/
8Vyln0wJZ4M1vAC7jHDTapcg4VDwmmn2/k3AIrYNF23eBwKRZPljwADkFQbWmYxIztM2zFj+y0jF
lGvjan6H/nZc4pqqGikb/F6LmLgSZKP6LB62kHJ9N8GWcBmxArv9BBV1oQT0K2U/m7GpNRF1xDdX
fgVVN4cmBeFY6idfXvBTCTxTh+pFyEfyEwcOZyCShD44XybemGmCV2ugXrfsJg1VLchIUvNSPaZl
cBYmykjBubjs9Rs3ERHcWDL/hLbwwXLcOCUBuaHnPvpiS32eeNEXIBnf2Alfxtnw+HHjuIwSJRQt
FWXgcxzbaH10sTtYWmlQbgtvSw71diOy5AkgPdPif/NB6aa5D5VvtPCJr32NBodREKGF6VfUMzL3
z6MuvNnqjprRdkaJEiWPlHuaiyqwZtLOncGf3A92vFigUMNWiUUNC5hOtY9iy5mXCRhpVl3EpeiZ
ysH5wYJohKGVhY/pOfMv39JBOwSIJuv2B3OutwaBdl8yrV0U
`protect end_protected
