--This example file is for demonstration purpose only. Users must not use this keyfile to encrypt their sources. 
--It is strongly recommonded that users create their own key file to use for encrypting their sources. 
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ZMKYtAygXY5kTNiIGmhLoloJg5cU4tnr2sksC7WS5wIvBC6IRbVL0QRLIWb/D6xf+nfgr6TnbZ9H
HYBGhJLGN/qPaJ/Qbmd3XXoXLEvvpPVmXNeN9/zIn9oFwE6TQzpVuLrDZN6EDg8u9IjknzefXtNw
Ez5mZ1nt+a3i4uEQJLfWDeWr6yjVgt+eJ5cXfoFER/ZKkfTJK6CSJ9amACUVum1EfEbm/XSxi/7b
NtZO5Hm+jGKyuekWdHm/iOpDMpiql7sU6JiJye3D4rglPhU4txjkkJ/o0v0/4CJKgKO+rEs38cEk
+cQBS1wGYUq+jwjZ2/NbwZMIDQjULHAowc+I3g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="zsPKQDeNzjurU+6Hv7cHb+3qXVWlcFexMYYy8SPWefI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21920)
`protect data_block
2dUIRhLHPP1uzo1SPshHCgYtsc2/7t99pCILR1mP3lh1i9dnWIOwG5iSP8CofenMaiU9Si0V5/sC
9sTiIhsZPfffxKv9swPHPMfHj4q/3xDKS/AXH8QDJ4zbhwJZfqEjEtaTECvC1Q08kwc9fO/fdYY9
k6M2PaiyPgNd/NjANbUrCX91BA3l8Q9yVpnHVysVcsS93vGEDsPDqRuNswj2MgPplFuJywLaPfhn
uhDdOkl8+zSZQZ8g+hri6uMiYhI0JuUwlD60X8JiUA+vi2+EU18g/yXnOkirpm/e0Lt0yn27Vwk9
HD7Nu6D52VnUqTfzFI0dvdQ6NB9wxUN+G1nxbVSX1mjwQmsVpiTVl2qt+VXZCgrfXAURHTlnQaJ6
fN+eGPMh1izRivHQuT/ceG3muVFRpxZgiPQwCjPIVhPokCeihmgmvEzM8tdwnQHOthJ0539GsP5+
FxEJ4PH56X762IM4NNDqUeO2xKGytHbNHhFHMOnMZYFmK6b0vMv7l+Gz8ha/GYQLZyIsQPKKXNwJ
4EWwIfjkfv016xrQxtJZVi6/CBSUex/DodBQPi69qf7xFAQVA7koA6bP7lagtPJygsR+TIn4GIrR
lpLOKuv3L4UqvbQqkZL7NGvYwF6MGZO712UER6l9sce/8mBzdQEbDLlo/bfCwEf+hKN1JaTmUPfp
P/8jo5Ab93/9qhgCgrl9xNYbkwaSjoNiXTCPGvNP1KA8uUW+SOuY0q/MLmbK9G0aczt1B/RDZBOO
vWcJA7bK13w0iMEaXn+qelan/ljAEwD1UAqdESqCaX0qZ3XPZf7Lnt2hf+SyeGpc2cnSXdVzXToo
HIWeTkMY/yzFUvAjYeicJNgJtFKcAvNTcAlmjxzuS93GGQV4grL7UBAKnp53/TxCUTyxXmtzyY5x
zWUf6wfTGWnJj7mlic8s1CweemR4LPWGyU96FDaUQXn0iPHG2SzvB2mmJpxbs8zUHI5gPlsgvmUM
bz0O1EPLM9e2+YLiI2sZJck3PcKBKGldfK8SX4dytI5CWcadR8OLSQDqOEUbb+iqjHcbzMODff5t
reI6+53TsnDWqAC85UOCDfwRTkXl4p19xkj2u9hQ2LGsKHn5jBBOnLgK9fwyep4SqXauC2yP/x6c
trzy6fln/dGc4uxaxM7WoIhKPHzPPhWG3e3t3LB5u7TH6VbzOvhssJ5nhcyrpKq6I+D0NOQh7dw6
GLRYSJkjkeuvtKLDzd5RPbzaDVSfb/Efmw43+8mXfBbm8se3aBhvT4KVYj9Tc3k//y/rBggYpGEV
iMXT9eBiE9Vv/YwBbDch5kktIdiR3D5KrweLR/gXNLmHUPwuRRn5cLso1s8IinlVNjdZjxtHymIy
9vU+tZMyqmfOK8VmXBrsV4fBITfz3/keQMjj/Jsa5+KzPLB1UQZJT+ZT79bV313SdZvt/J/QvjSo
7NlutCkEAiNtmNW+9/gTQYkHdyUn2MWK3h9r0cRT76/MvRNlggnD7QD0KBWB3b75/pV/SkalNgoc
Ie/Xr9nJV7letXRHNeeTsmCkF+hcxgCeFX/NNu0SuTUn0R87dAzoBaKw9q7hDAbWZVurf27XK5yc
bAkM90jDYoSYXTsoeGNxkANeA2+Er/tmqiMpmVJTpx1s3DGm1wfOsXQn8wI/YAE8e3oRQfI1ONUF
pdphgwv55unKNCOyt5vc1zhFTR++NG02DmmTZNtHdABGboU6ksCpKt2aZoxCqN5unD3HqXgwZsL6
qd8jNLEwcMm/1hnoMsntZv0hjaZxb8V5WErT81VUtNGtLif5I9BmCokjvGUdBPLxwe9ARfCSlLi3
V9yvaC5h0GWfatE4oTg5BQk4n+Yi4pDHiYQhGHXi2/WzYi837REiyOTrNpaEH1ZVHjamcm0fIUxI
kZtGEo2s5o6BEDw+mSr7meFwCrgPCQ31PIZjiRPGdxdX4Inwwl/pOcN+M4B2m1M067nwXL8WEn0b
G2m3VWIm0dWJjb3k2JJCFbMpBTmcvhmoO8wHdF8WChgP/chKjUYF+uzt+ciEu8TBupsaznV26GUQ
28tcFVPMJbYGhAsXnfWiXYVxoDrlUIzp58UEZN78MUGWxxzmYOMliom1BORp22SvRMkhWUSnbeYT
SjnhU2CEfFMSAMWvgl9GiuUwv21dFwmSVW+p6SK7acEJSK6Ax88HTXY3rHMU7Vug/X/2om84AZDq
goGq6o5P8A3/XFstLfXSGDMKbDa2wyddz3RZeFXluO1oAyKC1fGAI9GadTwf6aDZgoCIiE1WzNK5
BjMntAYMytDKV1jBSd6ll27iLoxR/acBi+CwaJ6uz5d1jNucP8jwrY1j1Pu8TAgmrwYwahgrdEOV
ztX6seaeiqCloy/0UnnLMbLj3kD1W0Z7rLdtj7MeuECJiGDH4IiKuT+Q9soRjyblTUKIBGi093w5
35+IQvnQAx2feK1K7BOJLVfESgF70H2G5lzt0VPqC1FiT8aFP0D04wJEElEyDZSbXszcFIfnpwSs
y5DcXZXr+AB6GRpLUBS2sgCdTZ6E4TKwaelUYuxF7B5Tg5RVbxaWEUTefnbmAsF5CJ/qUyxmIKma
lze++CwgllplPv2/5zC6ViF1ZQOLZEMM2YqRBle8pFEBCxRNFxSfXutbig8btBDJl/NV+3lo9Tgv
h7fHgkUi7fBUnXkCh4ttqZkw6kgnGjecf8j6u+5fOF9diIYNLX334S/gzxYA0me1UzO/k4CRYpI1
aQ/mn3cT3AbB2LQWA8AZ+jaATBGub51OJXCdQP6dS7IdkeyZRkFfzQRELCX/A5TWXO5avrg7susK
bJUFchgrnxa9oXByhEcihEqeNiHT/wiHB1LHOLzHK1q5pJ1K6wQ89Tkq74BDzV8jvZOex1HANDUD
zgzykA8CFkPNUYKCRPVEn6bi1nG1r0ymuLSSeCjFFZ2/DYIhBoyoc5ji71ql3PG/wzQH/bNWHOXv
WxZPTL3swo+aGDtT0viELK59JIKT5dpxXWDXpSbuwN+LwhYk012nDUW45kvysxYfp20dA/ofqtqs
Cuj8qOgbBNiBb7KCuTBnuPCnUFzJSOFuA4vLbG6wFt/sin7hJd7i66R6EbRNp1fBWMQZK4UYtbkT
YRB1mTDDUaWZ7x6nUmcvsQblEUAOqmN5b4hVeFP+Ot21AepBoth96qYNvSYKQLffyUoqk1Vl7H8n
D0HdaGpArtnCiYA3f0/GErExvrpBfVS+u/f2O7ZkyztmBt2FyHkcjj0IPyapZFczwgkB/+iwYqkL
E46NGDypXPwfFjCeW1d94lSSlhUXauit1dv3MnkXMHWdif9JvR1Bi6TL/iwhAobgXtWtb5ZKG5ty
tykNA0kU/qxrNC4wtP6fkNdigvebqiej7jx2Fi5H96FzA0sXrjhZwpFFa4lfpVaTXCjocPJuOtyR
t49JNhgm6oCup2TZMjwYM2KJg7QqSnuU9vhMLGK3b0O8+H+tXYQm+92/OvCP7poofBE+Ba8g1Hcf
KwVWtbihakyecAbX+ZnYnakYkDmw+pjdlxHfnTlAV64K0rPwnI2jclduAs/CgXHYFv+xcmvbpHbB
SYIIABSGhkuus61dSR5VM/u2F+f0oPRH0RBQa0Rek6NO6yX+v8h2UlbyxlpWnECFfK/1TVS2GprZ
VlC75sIjolBT/zJV3i1UAmgry60zSswUEC+bRWvcoSNpbrqORMux+6HWmclDcueEhIO6DTWuQe9g
VhkITao80GYqDdci+0FNVG6TRHTxWuO0THpsMXih1AOHIk3IQ+gTS5uXlJh8t13zo0CRxoaCshWy
O13gJ8PMp6+jye86oie+bGg6aB8QI+iQBpWKvjY9wcZRUayDLY7GIbVita7Mz5kxoMjg7Ou8wDg9
icAep0hVZEItlePZQ8NGkYodRmGGwhCHuP5I7QNJFWxhYEzPcqBxz5Mu65oIc6SbYmEk4QVpk2as
aFSmy38pPRL/FbE7abenxZyhmlWYUWfPn14vttksb58gCdaEj8pRnVPPJ1NxokgAByk3E3ND8Cpf
zWtJMcqiUrwJb8QmRfRlcbXtU5/gVwHWeDqTJgQgwOqr+q1fTrEk06KW/V/JUrsBVsMAPcNcq14b
xkRvfFz0+JTzOrCya43I2840uc93JcyaIjxR4OnBNY/Mf0xMAfVhnM9Z9hUtuCqMxrIAuT8Sxmtr
ihQTyNz7EVKiOCWkDxdFsiz3kCHyKoSkke5MvVj4i1duQJyg/kqfahgAtc7EFRLatrwdDj71nqqg
LNYvuqYFR1gdbFxByuq0LuiA2TF068f4LOacmr+FZhQdIh3RZbUqK+D2H7jmUGdR+cqJzEKgjg6M
7lx6swqACDLSqgsXgWIqQlpM5cqidtuZ/UFTHGWhehAMzPlN/Wf/W7ypDRd+5bs5Jh6fef8njveP
P5XpfVWpiJ8pneKa69++9a0yadTMjufUTJxmFXJuo6caEDYkSHrgSlq4e5SNG4dF09qV0ArKoppn
YSm+xTpJ6wSqTzGVl3EJAIBgXDPUkzVqH0SRgSpAQDQ3u7pUwYj1dbqx3011W8DH9o5j5mWoyWMp
otNeuEihrmr2vTl1AVbzn/yGkpi8nRx0/nAmvYCbkj+7Z3jvu+boh2N/ZNDllU4NrurRuyXATdDf
Bk+rUnbv0NQzeQLy4IoQ9qS7BAWBLgnIJM2PnJ161OwbRnrFhpWFsvwpjBZK4+abjW2GLXgia2mr
cy+WlBjyWjAle0v2bfLKy4nMUYKjM7gGZcB4JtEalnfY7DuNhuth+V3K+/wN9MpEMK9LKi9T0jq+
/y70pOqzq9JaSEU59V+dnZ+ym869isqqp9I8W6YwSSEDymf9taFdCWnhfuCHQL5oDOqU5kOSmu5p
613Lj1phpXzoMM0RHDrsgWvGGt9zbmeZvWbEvS56KHGy4fkJgC4tkBifcVYCbug6K3dThJAK4MMf
Z4zpjcXTvzz8Vblu6ALn08DDGSMofOseM8MO+QSEXAjpe5V+jOF+G6/xZTOlR9q6rclVCxzRKY77
SgLg/fvzNuNQQfYghrv7X8pDGCpMGdFNN2qppTN9gINzL7CqQ1JnLGVTr4rBab28lfRR5EIKInZE
aD9Xqn/Umkkh8OqMSM1lJ5nDS7kN8O6i3X5O9qWP57WrG0US6RhiGo4rAE8ncJpUd/pAgJ8GVfUQ
HTFK7Ql4lP9kKFcW9CFKVeJAUtE6b/K+L3gQbO1DLdz+as84dAPu+EAkubVXnhVg4bzOZhQJKjyY
FBRK2JHcpKQk+FCb3Cq6NsIJ4xFvJenjgDZOt0FgSehIKVwaTK6ecImFANUGITPXhkGbI61qvx1L
CsOvPGniQ5A5trFnqK3C14TvaX8QC3SC8G4d8UjSlAtjXm/nWau9JkWaHvEvejm/RmxZtNC8Rh68
GpI7+z+NUNketv2AjQ7yUASGG0VwN7nz9yZubGhtFlKNPjZy/5fv7NE7nFxQEOqigStacFooncod
iA1JvPVYIGOTWzoGxUbg86XHJM4YzDTpQNjrbddZN8tUwfi5/JhJ0IsZG9rDhEmw6hZ9ZyYm2ifM
/93RS+NYhhQnpemy++HOuFD3bJ86btPNb2qHL+ISMrFmlekQAxr5yeiTtvYHhQpwA/fGldS2sjB1
Od9SqTArjil/wU9IJJl1OM6mGIou3sM8ZbAS3UpwWCT6tOJ43KVUGJtCDfcMNhgptg5jep0hFJhM
VMjNXHmyI4xcYaf9dfWRo9ssGo+bbxjxdRhEmAV6wQ7QkxOTwixth6C51isM29p2idL7VVbNOrsP
dQrQ2d+03cuAKr3+yqCv3uKziUJvt5nxFsf1ShWFWcoJqE4NfVRUh0s2yuq8HaXrOwIPcBT8kBuv
nrH+m0Vvmkr3YTC5PoYAeqbJX6OPWZMEE7UeOr99slcjqc2HiITuQq68ie1efGHrugjnMeD5U8Ga
dvRCRP7t/mFuYyl0dT01u8XyLnyR+FLImNZisLVn2WWdA0RB8We9EzaOIsABXzFN/GBz/tKMKo1q
lLt9I8ZCjrBB82xyCa6/3ndRPRllCXlz8RgpP10kptyyw0MnfA1oGXRRbI4DZeEFKTERulwxbDiM
SDb5LJq6iaKcH3iTOaHi9LpTwpe08vnwEMN5lfjY60zwYuRkDJ0Ezh75Cls5nROlZZAj4Ue4hX9T
sDkYKoz3mERt9LPtpNeWwu1FEB4UZ41Ognl87UJ1637Gpry6KAmqzgvqL+VNG8KGxOY4QFYa9uGN
zwv/YD7nBRMFTCmhRUbS1+ZyNt8RvTe+zBWACAjokw50TTbbToz/ZqpwhOifDp7Wu+u6McsP4Nya
3BMDFCewiAAA0xgFShFxkMbwahVKwnwj6D75WaS+N81pJuww8qcBbnMDqJ5grIRMWx9fhespa6aR
0kXGk1ii39PErtmUvDGr1indUnJ88mSgygNN5CcQcuaGUiBNY3HgUfuFwXcw+eWPjjfKffNaGlNl
8VdojAFxWtMCIIR+pseYtT3fz19ztiP7PDydyUCDNnQRpuc7S208LOlFnYBZdwv4z3EV1IQyYbJC
nJMuWnQCUbPdCiF1vnGAylPj9U4CYSSkp7IS94WRb4IycfGKkygC/ZEzTIOh/6f24S4SLLlqOWtL
AzN1AmhFmOXPMGEy3fLxH0mQkd3ms0yH+hPNSaQ4kWyxWbma3pi3adiULsDOuApnOCMsa3z7UKjc
khoPfp5d4j8S/r10AS9V84Ec4ZHSrJFaXoGNiYXX+yXEBMbM9n17wJb+Ro6kM3N+q3DIU/EbeeJc
0Yv4vu+ZlWAVKRxatfv5R6ffOXUJic14+p5WMPiXkqWWGMWwJK1te214/2o9/LsYNOHWkId4oAp4
AbDNSdWQFc560DaU60M/ttkMh/GqclwjLn1JuUdszGwNU8aKdMRgco5NVdG7EsLO/2TADAQcQo4D
LDkrmNh8r3YimatTE+eYom6K8HXo+rsEGV141kAe+MbJbaxVdu/on2attrRvuXo2GHDNUjJ9W7Qe
Iqwf+yZ69g42GclUf0f0uQnDacazFe3M+C2gySiAKPylWSCFSOSrSe+0QHH0P2QI/+3AkN3qq3Px
EIcN3f8pSEdJ5SMgB9FkgnmOBOz4yo1WD9yFhau7lUWuf5r/SlsdPG1k4TLzwNkDmii+yJsMQ/DT
Ioy0hE+wabpqsVAFa8WVoeKZ47xpzGzveDyYfZmDrnTdXv3KCfynxe+QjtqWamkqTFlcZgGTwOMD
MJil+ElpTBZBbUuFtTweJM5/kZ8wHnbP5ySLvdIX/HZcgDT/a55CrlRUS3kJLncuCUWJwOpISKxB
hHjLQV6oRHJ+o2r7ggFAApUVkg7XckvPNAKHDmNh3iOkC9k2NlitSe/CK1N+nzjeVtRGq7zjx0Nh
iD1DqSMs/dvlJVpc9NW+wPr6lXUTACkIwTu5kqCfQ+NvZw8L55le0f8Fjrj6bYBRyPUtMLVN/Wrb
ja3LEWR55/Dn40hxi9SxcwurhmiSECP3oY5F4IEx/fSg24nGHsJLmF836D4wy0xwH16bojYxMKYU
Be8up71Bj4G8JgMcviA6JAMjzcgCLAA54msCOV5iqnQJDA8GJlzd23BEtrx397btiwFAGLdip/YJ
2SOmJGnN03jomA3DcozCzYYXuJvktFz4c/e9RKD3NZ5KoOctgxwAwY56wPfRyWTb2LUNBGUpA90y
9TJKzgWjW3Jze7pDQtAE92LUBSgttm289XZQHjfBFvB80fZLKrozIGtVzaUk+sC3tplVjgm9Vv/3
8W8hwl1BnVGWFF7/7e36EGlYvDW3SttSRW2J6xiYxk/uBpVDUJoy/GxfWlhbRo1i/7NCuFJeeUlk
6AA8eEVMfGNQLp/5+3uh5RnfIvdVE8x8Oo5awCahB7eGQxIwnc10utN615cptfidjsO9BfIRz+mT
77q8YNEfBSBbB8VTl3v9AymkDQHNbX8pN9u+9RWngZ6/svq3GlPImHKXuA87BxNoMmpNBWujRign
Lr5bUsHtmnlg+OFXlEF4TLCSwANZljNW56w2KwCU1WVBmFJs9PdXdB66Qx0clmi0Yl+x26f/ZR5x
ykSzLmwnI7qhHNfVbHMBeUsY6E/cEEgs2jNks4vQbB3EjwfVK7VGLiHqMwg+F8ye4JB0edy7ba5T
pNXgeiLSGNT2X8CrXiqVQkKmFNmHLJIlpUreTvm4JPf1oUQ5l5kX80nSFK2Exij83xzWg/w9k+Vh
ubqmZBG47yXP38NCah3yskhO0QzpT7dYgjmYpx+RWD2IdqrFNdcYJQxkVb5BKb5TOHYMWpoUEdag
JTfrUumM5WiLvcVj/P88qDlg429NsN0dvQIp/2KGNJ9fLbr9LmacbFoHrD3UxRiwF4znFKPHHvRX
lMkEiOI2itKu0G5jahAKAYdqbx6PgYBEAkzYqHh5j13ZxOIqe3nXbRluIBPgjl/lpA+/sJO2CWaz
ZLpfjF1AO3JQKcC1KO1yBfDLydMTcQmLBhb0r7vdxe2iGjeagGgpiuAivjVdlEmwxgy3EOsMG3QD
UHtkhmGiOaOTSPHqonhKomEwnY8LeAVYDECgHLAmuXIBSWREnaaEauxSOZUDlYIM5p5bABVe70TQ
zHZgwvJ3yT0htEwSXm0KQDlhed6eoildBMv+/1ig56FUmSs53RgJLIYuYJMoS74ruSDNbk/Iyku8
ySpgGco17eqUnIMPgkmoaXndGEVWqzgCv6yV+HsRLlfAcR6dHsB96yfWZLuXCmiCgCHt7+PiZIWG
m2RFVP8fTT/ehmRKvKseiHb3ilZ7ZMP6mh2kpZs9U9TfoBJqZ5OFdWGIea90HpHiYAxr7dYOqDvk
3wKXYXg6dOzp1wAn25yxvDzyYG0FlqIecg018AZyR6HthG5dL1njupsYN6aYsxEJkNkWlOFe6uh5
AQwJpxPEM9KWvABkXmlW+x3MRCUm+Y9PvCODzReG/AXwTdbabM2JVLn0hTBt5aImPL7WPCZkvJed
XJh9HxDVksTYkig6VyJTwdQ6BjAMkW2MeSyQ1pEl5vNWEHKA89CwfaG1HAOCBDhI+yXkS75VH7fR
wUqhcO3R3wyMlDkHID513q4MX/qY/91u1P01JjpnagMcSP0eHcTQSej+FpkzSkBM7idA5PTm3j5P
vzMqXhDw+ZfOSenrbaFsNEO45NU9M25gEnrVdRZ0ZZHqhRGHCiYFh0Hj2zxF/XO+hlTHnBEOD3b+
Elw4sUFlWERqrBcpXUj95dZwM2NC7ere8demqSYN8pcqlFabV1goQi4WdQY6IHNWR122t0ohVvqC
UsGl0wYjP4k4j685dK5aFlC3/Q85CGvfjaKP+OuCxlsj6OU1h7EQ6oaAluxScj9ub2GiV7q9FXXx
u9E0Y7h21n96IejSDTTOqyvknzM62zPd6ZsDE45a1k+qc0PHurJe+JRAZVUz4sdNsiU29IGpFMzi
baeAb+aEEB+z8lZkuvVf5+5czec+98I9rBk/AUJsutM0oxysrLb1nWDPhUcMO4Wp71XYYD9r7i1l
QQZjFHKoKJeFRZJjNk/RWSopPXH76wzbtjhJPY8DVaymvKgpHLqzyJMv3z7kokjS4hrh010x7XLu
7c59kKRs4Kt4xf6Z6mCB2MoGJza2saEZJxa18pjqkk6TDKpTYhPTLl6cekAv8JEhMSVJsEkEwmOo
X24TNptfNLQvuR4CvjVGYRHjPakAYadrSWnTE81rp0i8sUXmDjGIDIPB+uHFltjbW6I6oNl+JHm1
rbvUePPMrP9UBhGHJmlxPzHa5NoxP5gD7SHSdG6Yqsq8DQNNp+ZKlA6bpWhtqqCpxFknxrwp5Kp2
jPZHBJomxfDSrUhqUpYl/TYm9Rp7ATepW0jt0AG7REN3/ugsRSHl/TqInXGMOpvRndzjVVz9eLci
dFQFdsMyERwX93o6fgRHEWvnTW7+vT+HwkQRy5CvxOorCX4wdjNjfbo6HNMN2pwCWmYMzumu1uU+
Xr4e89eX1cwzu+EnHa5Ie+S1Bwmj8LD6lzalPeXMPMtIXCQTk3I39u2JbWGEzeB6qew2QTQR0Mx6
o5RvlAIb7YpIqs2GQqGUPN+U2N78xqXo5hJ1N5UDbbul80E9OHJpVWzvxf6hVJIKWJoooTVRI1PF
Q+Ll7zBht6xlYZtFr8WcL9fFEWeFU+a7VIrRrqMdbhF/ZNEHh0GLkp6FEk/k/ILOl2WZD1FyeXzi
OCRNr+DtcgffjEL6mKwZwKFMiP3V9OOP/550gDvfOBmJSV7oNntJzikCSMIVH4jdG4fM6+kY5b73
sB02ukbzrX2SYAI1Tls6qaTcdiqL8GvuvRpnxCjepvuqilpjN4mAt6vBO0QfzRm9+RQxraaonehL
q+2ijwDTnQX6zaKDE1TNnNxBOZYkkYgvLcua739bNGUTLtrvuciVguxkOlH8VtXCvQRfjB2b785y
dq1Sb29s7gsPZbYYnCzqfqtlbORSnVNt9pTWPbHWvpatH9oMN46mDqWr5ONb3Nwqt0oG03q3a/Mj
DONKM4ppypxlpuBBnQmD1YDqflLXjcgDcrhhDwqOF7vRO7qx4mE7KGwM6HhdC8tAsMc3yYbjU3EJ
tqLZ9fgaWkiqqpcfPoEk4R33Ske2+z37x0DRSxjjmGQRcsa30xe6SzKUGHsMXwOtiwgJVCWY6gXk
Tgwrkrkq9CD9xbThw+mOnfvxL+KidOLKYVng6Q8mKGuNYo8MdafoogUhMoSAxqhR+0+X50DZiWLv
3cdzSDztDQW1/INXCK7WBpWVldWRw88TriGT9tst3xOa1uqF/z9BCvbbsWbsun/DUXemn1WHpo0Z
IN0rQdhLP7iFAv5xgZRbd6jwUo+hajsMXVH86R2hEV/fXhL26TNFANeXG4ZcPKiSN8j+Ee4ShYIA
t0YfG/EIGJteKxygp2HHipqzO3c02nVp/rHatVXxHwgWge7hrv3EVmJxOXUw4MjitcPbgA1eHYyx
6pY8G7baVPhcfQfErd8Fcnn5m9WtzQa6aXep55zrpCyQtkv0lR+mRV4yp0ob4vmxYss776eAJPGh
/dAelMX8OruwbiWvAYpW/aEay/4Ru/K2nBtAVFEmB7VordLDsrJtmk/JITUuYmj+UhmkjAqyhHQL
9r257pRpJgyDc1msa3Y3QrGtJPDYqoh8LpcIGrI+FTt+F+Nv+J7Z7xi4p3Sy9CWSZ3ETE5PNeP2A
1ElyV5o5zaHWxqnNXnIz0L7UdIZgryoWF5xYW7HBPBvD6n7gn6ysewu3VQmqyR31Pl2/vjKX0lJT
exnmUcij9K7nxaJjyFDVF1UJ+J0lBeeTkQdkCvEYZ5fbxma4IS8iuNpng4qZaUHHpum22I4kaOWx
QIJGZ003g3aZJ25uu+/siSaa7e+v+xAvYehJhrcI1WKjpTIeIAdAAVXmivfpt8x1Z0Les3oMMdg4
Qe/OAdPjgdD3gvm73spCdI+dsd2V364ksFDsHJMZRMvPq/bBdjba6KUlsEgNtjP3M0cDkcY9OE78
nLmBg7bOv7hJVH0d9JjEVPVNMnBzziM9DA3Ox81I7Lb+Zoskm1OMu87vXCJKQmPMbIO2KNsEajdA
RHLYAIaS6miA+PzM3yunTiZ0AevUdOSVYHoa3KsG/jMGYD2dGMvkyknqjXrpwML67PpDv8kDK8S5
bE3f6faYkNBrlAjwIpXeyURu1ogyTUpuVVz8zZ7zmFTvrFX2GIDptDW99fgsE+CliBE6cb1mO6J2
s95pS4HmDgwXSRZ019IK+0rV2UQ+hHAkXKteD32iQZQs72XIpjRx8RWp49Fy3JqsfX9qp+3Dgm7R
jFS/4ZjzG7pahwgftxXehjgqyTQV8ffpsNhmZsT+zIg8cOmMAhkCGNY6kCcVu10Wrm8WuZyQh8Iv
nz4OTNKF5LzWD38PMgNr6CdVrn8i7wTZrifGWBx5iGJkwt9QR7cyPP8q8tmlS0gL4LPplG+ztuMo
mnjHUirQK/VJ1M4lqMs/N24Iay7dfG/S1MXxKUVsXYLKhTYWb9brvQhTYq5sS3TB9sxB0cksAB/E
t6MKpfTr4Pey/oVjZYddsCyoLOjmIyCNmSrMBY1ePujeckDWEWUbNTURHDy5XdlBoNGId0JFWfRj
N+g3sAJykrVcoGjOvKV5xeZbaC0zH6+6fLfl/tvPcjkg0lGlR9cr3FNnmSRODiImgR/4B1JKhDy2
7G5MdEpvEPTQViJrb6S/mcmTEGJEGcoGLa3q7+sVPflcJYaLAi5SIDaSH+rUHdq/amwXl94hOZQp
FTGVGu8UiyquMRZ0kM5h+4bKe8MX5/jk2+DQwZedyMmN2kxsRWpRA3a8z/+XzCCg9Ya4RDXQXqvH
Ye+UVlrIwcImQcmR9QyLn2mhMvOTbUXJaVLaZt8c5Mg12bmJM/bDwN2vkfFKuhKWd9+CH68pjpI1
t6eTuIKX4D7gpFAum6LGrhpmHcF3KXILoJqQTaRVhtSkrRFJBKQR0bPVpW26O0RUN56yddQCKnUB
eEeD6GPQyRw59kHV+t5tXUetNVq/VTEn7D4/BmhQCtL5A3WBxfF1HqLJnYZ7jNO/t/VbORCe5hT4
5yfIlsGbPeiLbE48hqr6I8GiNqO3vUBEdJAVuoIITRxuWv1128I5viWSc9KDsM5DfxjcsbOCOkZg
Jvtt8smuejoOURxparw5wAv6UMFe8QH+l1WrLbvDMerQ1RnE6XUmQp2zWASBZoe0ytHvs4s9aLRM
deSPbXEJFs0ZanwTwDAdFqbcPfg/84VGiyG3zFBpUGNMoEy1yjt2II60/l0MeRyXWuVtyaiz8Fu/
9AQoZwHf8jjig8KrPreI0Db7UBAOzg27aN/cgJOYywdGgD3ztTifLmvD6Is13BXfhZZH/MDKSOZS
9Pbw09P3tYo53lkHKhJBf09noZrDfx5xlRQRfT0tYm0WaeF9l7Z28x5AwYRrCU/J7+Svj+puOaSD
FDgw/lqsQBmyzXrpWqdxbrTtEi/vkptWGV9QZeuyTjtH6CkAhMbV3Af4CfXyAskBTyluRe/zJ4cS
FzEgTWdvmBagClBIoh/XS1JEm7grzuVurIGdo8kX4ERD6PL4LL0u6PRPzSsDWNbeVfv0MnZqSSvt
1qsHp4F457iSBoOndKvtVexAGb9mZlXQNyC/a931VUXdPuz0dAk1n4k0qGsqruBG2ftTSZU3zPIZ
jK/QfR4UPDZf8LRF3GQJUWkVhV1LqRcHmaM5FV7t+VZ7/9mPPv78BCBS/bgwTnNa+M9mdW7RmoD/
h2KN14s1ocbeHoBGy1Ggyn5y0inijBZ8/lmRN0A6AMKLf70xICRkChi9CJtXgX8YB9sk2EAIAMDr
FdTUAtQOfJvdxpjwU9kG9eWqojyXRmVEvaWcfDEAG5xcEsdG+9Z7R5XdJnTLDMQxsu+Qe2yYHtSl
Of7xurnDm1rmwKVs/+5TYxVYCaaCn4nm2wmP6Y2ZPvcea9SfMg5EfTKzbEvahUdo7VnP4SDIzBtc
TwbJhkGkTvUzVpZCONqF/rNNQ+XBakiylOGlaWuU5bUH0ob4roG/T69VWZqf5i8R722GPiCe8iEY
hWwL6FoK4UhY4/YhfsRTj1HlqSh5fvlM34eV3KuOEmlmxr9UhwBRFXWP1ByNwjXxvKEV7jyJB8sG
W1bPwG+sm/9mwUkVLiiXnvUyIijOw4M4Qgt+bQNr+wGrQgB15DPMXiua0DHnWlyyMbng8G5pvowB
nwyLxlBh4aR2z29eXqNchpy2XeuSr0l+6Qzvwq+KAHu5hyqjimXsLX89WlOEsDcnKCdVGoIqvf6+
m9qYVMOcFUEdMbL2k7BNtvZqOAGSSaBkStBPOO4SSyxUgZrjm6wDv88w3T6Lot9SxP0ZwE4GNKDa
cq4CrYttfkswNb3UbfWINl2iq0zfHpo2bRmL4zSQ4VZk2V3/kJPlpWHCWLDhGUB5yyZGUZpjr4hs
lefANEqX4MkIH5RvxyDlpTgTvQU8ESaYllaYuGwp0SpulGgs3jVLRUbORA52zVLfAxDodZy5Lkky
gt7Nd+AQEAhWCOpQSouCx+fW7+9BTM+sZRMuYwZ3b7lalbcIWMFqw9C8EjtEOwJy7mfk+t5rZhos
7raJqunt4LGAWNUMnjnfxStk6+ieqE12fssiKj9bI/GtIUAegbnnNRV/rDtYdGYF5QZYU1ucJRTR
6uW6P+ok9BAN8wHCP94N6JXizEfl5MDvMvBE6APp/vnQ4G+fRwAGodYaH1WURh5VXmBxDbHRVav3
5iaqD/GAdEd7X9D0Ex8knwAFaAkZwXXAEkg81r/69iICG9OtJOzv+zOlcftXu7HUgUN3/G1mb5Be
k5LOEokhsGV5CK24fd73f60AUKA3jDN2+n9S0ql28gq2ciIXxUK6oKSb3iXHz9wTiFuEyMrMPxfD
eIwAQ+199eRWpAjXN6SE86HuVBWMfHjFzAXAGFu1ZwflleF6biEKDj+4j5iCf89i4LwTA8ZJYhUK
9+Y5mKQOyZRJAFc44JoZRRPJtXfKNvW/dgg8EpzzjZ+l5J1xe6c3IYfqikBm2kHdtZ/ZPkDXWpgt
YVkxn3+eQhaDBddQ4mtij5XEOjllk6vRGr7bQabv7IRHUdO+aRXWVQmyaOYcXDvqYJCoJpv9Gq5D
uAwUgXwadTj61SyyaZEqyB0pNi2D15y+IU/mwD+ltjxRfskVNSh+1hluiNzmWRQ8f07m90VkOex7
pGEnKS+m8MTnR0HrMjwd3WCg47zX4hhTsPC1mFQisKWRUuN9oZ1lBosuZLW1YsF6YgKYE6hc+TJY
WsVH3G32wr4maG23qjWmtsELio1Uda7yGlYh4pYwcSM9LYYeDhuAXC/z0+9qKizGVF6meJnCLNoX
TUtRf/1Dugb/TaW/0tSwsCjuFs7CxoybbBxLjos2RqclxNsr0qgNKmONdk7kCFa5eAzbPrLBM9hB
kZ1hKTYpUra5mG8npbEsq9X1Iv1AYqR7Y9ZmpQWJu5j1W0aTxK/sIpF3O6rYE1+XxOXsoqkshOfK
GwbupyDZIrzrgg3Mdt8SUmL6xxiFUNgxIPPbPng3xt4poUN3ft0y4HEzoELR7nwFcCzAx6Lrizuv
jGJkr6CFOLFt9nJSLVaqh4zR6AJGRZTPI+ldJZcW9vsQXa+YvUnbjASLyE5xb9Yav7VUNt4QYnih
+7nJQTRFIpullOXG7ENtG1HiWaxJ9GyWfS0nVj9IrsPXdB06ZEMCl5oZDDsm2z0y9wtse+aRyj/H
FoV7Lv0Gx/3ktL2CuSN0XPKRJYcLk/u3SSrK8UPX9vkw7Zv4uRgN3CEOCUkA2BW7j2bOCZUrMqfM
qz4m4obLIrRDZiZT4lSe6a1Nd9/N+/fo56GvtPYp6Igwi++bFezQyorlphNv6NCmyx+5uOJyjihV
sr7nhCZacBV0LDE3xjAC0L/NwAKxN7/nBTpyxAsgk8FmS8SdJx8e/Lw72g006bLk+GVOf3dRoGVS
HqIz03h/mvBf8dzVvJXslJnJPfXH4plKbm/5eL78qRNd+oZ1gMUhpnbNxzBe3C6qdpKpJySY3xiE
azwVuJAh4Bq9sjJtS/DWalogHmv5fOHWWCVZpdNmoGvGRUa+oB18bzOjc9lNkt7knG9ljc2y1I+w
QKWqhG1h67uK8d/MejbFWznRFBseJg7S9Ogt9sk3HExpontimvHqSlV8CY24opck95SqD77GWLlS
kYefg3Eve/0vDED9awMtr76fx5+AcDQ8tZ1bYWRhurjwVd1GVoyn09HnKru/tV0KPBAHTKiARm6r
UWbZDwZTIe7unflWqB4/2mkRmeKdPpobX7yJtIznC9I1mDRCHCl7ETKx+E2K4wFSrno8ruWa2i/X
iwHKmpj+qolPLgMmbjFUxG40VjeOoUPj3CShpnGsbXvd9w4ExB2VOgenxqsik6Td48qEsw+YZWy/
W0o/ejy4fPUX0SaKjgGVu5OIjfik6C2zfdxVGow3iXfTk66judRiFrngTGlaCHy1Dm1LgdvZWgES
OlbfaH5Eb9Cr+zMN+HergzFDGXqA/h2gd6QcriXFXZ8rwsAYmcMWdbyQhKkNj2ndddqv+F3NUdpi
yjjy/AKwvUmtoMzZGIU7xYf9jktslqPm6hRxL8UOa9el3YCbxZCgPcCxC+DkVUQouswKHYBllTvI
G9EDE/Wgw6McjNijdqovJ+zL1pEw9AKQmTh14og3b071Ds6FcW3fJa2pzp10QTXm9apWqYKXbR3X
AO6DYpMoqhOKMnqS++tNsNGwppLk2uOs7XQpzZWVMKSI6zdv13ZfbInWqmMxslRJ7ai4joArhuC1
YwTZLKm/bGUhnTHppf/+OPkfUuy2kVswuOMDNHSXU5I7n8wWVvtEUNuI+dGTBDS6u4fxfpWHuDUq
GqYztByTefciuZpFA2PnYqjvDX7tziolAn2yWqYBQ/zz3eJoZr3AFWF7nmTI36eiC20vobkf3lI7
bx3ScKXtQscyFa3+8LYpsoPatzYweOGivF7FxzBR9Bh7YilZjKXro2ic7/mpHuHzzmC8YKAN5G1O
TH6kGveTbYdmhMewCiwuMiepyPvoFqQaMjFoUFxSw6jF32peUu5YgBVXkfJaduriauPfGjji+NlP
GaiJDvh8EwYSJq0wTjWb9YQSJzRh05p7yEWFn/Yd3DequcRoWTlFHt41/XOSIXzJhCkzv2UMQhFW
B3t0xyECBZ2kj5Ejo6AYQLJpgnRLvR6h0yPcFUbkF+jwv8i4tkBUaWsLtKDLjbWQW8H/qm6bC6b+
XZaKh49STswNtuOXLPfu6lrtcJDTjl5or+QCiFa+I8B9klZKe+DiangvjrtuOah7kJV71966isY8
K5FJ3JIyr0ECFK1QlbzCxRwNOFjKCuUa0Th81BQW9mEoN4/Yo1DP9umYEYOaUrYWXU+JvAT50X3P
Txq2CmLwXY8mIOWXml/ROk/k6761Lk0cg/fj26rnfRfPxQn4BQ7F62ldh3mR8AdSuMj8BHDR3QsD
7HxqgzF3J2LLGJuES4WEO32ir0fi46VuqZQbTeKoFNlRD6Uc6pZrFGXinCkBdU+MvPkquCIJgprG
fMNijVTppJgnALMq7DQcEpw3Ho7UGUpLPvzXlNIxanOmBXHDY8cvAXBFlpHKd8T0/hhkk+qzI33B
gfmxv0vz0AAUKx5hAQERVlxVba44p4AgkzIcGCOsCN2qtyBDb1iHzf9RHe/nDqLGQLi5gt8nz7hR
96Aknnja7bkc2KWlGgiZuBH/wQq7uO7CtPuFPqC2OMuAxzlRP7Uj3ZDSI0EW6CXKXAuX/1seZ0gu
hA0TXJNUkg9v5+Hcx/KxzkJf/7EerjOQDJDDBBL5oMY11VV9obtd7BiH9wffPBmA2loUbjWXMs11
wZqE+qEGSpukRzsvnMZailW+gVNbJgJ2nEApsKHQOYumrzK7BvRRWhG/aBcD28chOtkkF7lyYr1X
od0Z+LOCGw7JTGko3hiPlrRzfukCtsW7DCiSuBrOxRyO59FYVqHDgzTMeiZsco8vy0xcJiErJOl8
950brVrNM0Egvf1hZbzo7vGPEztgvKh/d8skMaKkLWFU4z0nONsBNUx5YFgQ6cGLMpwJtxP3fZaC
E8oeiShOii75X04LyI9iD9USEsupp/yrnDKHd/RAZPatORLIGPha4C0vFGNeVecqFQrWBcd0OhXx
QKx2TZ3rtAjby6/fX2IzitYUQmhSGA4tQL7oFNuTAd4S4M+1e+OPGrBW2l+P3tkop9o8V89u72nL
X8ijCGWmIsmtLnEC/So5DaPfhWkTK87gZ+7XWkk8GT197G/p+naO4cyTVloFXZdjMsvZbGSURv+S
+LT66oMUm4rxDqDasCO7xhB5YJA+Vox4TKwzHHHinFWBsoPWzl60uJASLd/NXmE9aApHcE2T2vlh
98bMruVB6I8xqADTewJTE+FKw2rPTbZ1eME7dmuPDCI/fPDRhK1Zfr321Sut949Ga/YZ9aINCJZZ
Vpq1w3XIFFCc7TsBJ7TpV5cZ8CXKbXDfgMDvO37ALPmkWaBaaN+MV71haT+sbBun0GRQsOIbvsJk
LoqyHQLOeuR4sm8sA5zrTlXO9+Dr3DDOguXkbls6Th6WMezWtkDAJ/q6+ZLpova1LWWwx6XkWdpC
IHxtv7Z9Fx5UCp+yi0bpUZ0xC4b7kQOCHlNxrqHXq1JyckN3RoZ9Wx4qCTk8eJ8wLWvQysrXHKbE
NZ3yNYL4lgaaKI/ddVj0XWntec3kU1lk5bjiGpQC/qD4ux+aN3cf77aggm9ZNiNK7AyyX0GTYWOp
S9JUIe9rIDTA+iX8VNAxVCy0wqbVmD9kfzWTd84gNij/phCQdJbidd7N94I522F/dbqdqrQ+P6kp
/qDhLMXuZQkFvXLxIfRI4qjWKNE63YeeOMTj58Lqoo3cQwMT7S1qN+4e4cmVpmpCJ89RJuSltuqI
d509SOFWDeVWYciQYb5W84Jq6rn3ALR9KZvlqbDQhfGmLp4m5k/R2MJn12e4jNpJHb2VtgzssUXy
GReJtfJZljtSrd0p+G5DW0AC6c+AkBXu83F7yXLqm3wQzI32anhqVvb2+aSYv0IJqnooRKNRiimr
bSm10GQcYmE9vY9tXb+P2Zvc94yvQgcN11kIhC2Eu/cRIOVdIXjMw67ENAq5ksYox9yy96hlbvmQ
2jWXK/NufgpoKoh6JJKDl6G8fb/DxYKqW9aWcpDIhN8U9H7zIHfE0sp+iFrI1L1r1CRHP7rpEol8
vXyUHKnb3sDchAk+K18ntz2fVy0OSMY9nWqDPYftACNoLWFUq/hD/cUl7hKRnlkd957TYjahHi24
MrKhS+T+YuPbOH9jdC8MhEbJyQVtxRYs5+/MDkrwulJYcUXrnLGBhc4L6LUZoekttgI0zgtjPdao
Z71W3hTvKorD3rfS9Pe1wY8JYyUa4HpGuhGjKwjE0rnm2W3qmap0H89HdN8+nlu77PocnEPpViqN
3sER5aL2uAUWNrJSyePI+TRxHHNIcKGfdjfOGTJSCIjuI7iaYEQvb7fK+iT+n7A4/CODXWg/BlWP
3WtG8wlHzsRxTnyajujJCZBw//SNzCuQckZfhiqzEljOPBRTNYAkb9hJouhRv5dAUWwZLJ2kLexB
j7ibFPjD4FKIMPcfDECgIU7Dvb8RWsX+qCeWvrijSC4NyZJ4fEUjLLENoVKRx++ZIvGvdFGQsP6i
CAlxgo33ALOv8HUt/CIJKIu5tuDdWandF3zBGB0vgWD6/3+oRGR7kehN8cckg42uf7PN0myVworH
rzDucYklKGktU6ETS7PBrSsICI2zddGcCDdU9e5JxIfznk3nSx/vQm7bXspmrx5PV3ay4Y6RkzLO
dvDAMKWBQinbPTJ31nROKEluIpmPEOK3LUgTjeXTdcIw12pWLmbjgs0LGR+NTJF47I33eW1sjCVw
eNvc4jhbHbdZq4xhqlxniTta6DZx6IU/XyQrbJLS1JwkdBh/7Dsugr2JhhdtcU3QFU8lzDL5NoTv
WJhMZb79lio6u1vlLP9B4bjE4h18iq6hDcElokj+okuQtZuRZ5Ny12S1NWaOOo64ECyqUlX32mIX
JOwVIBj5WseKftdp7GvzVVOVa6N3uATvWnSgiJOG8Ku/j/ql0lC5cFjUK3SRKYqs9Zo/URuRbMgO
nVuJTW+3W0xzW4w8+zx3Oy2nB4PmDM1ujy3ST6jNmwuCek/Xg7YVnxzGXeaGGPvEkBegJVHVQlLg
JLZ5IbDfZ/wEfQ7XUWON5vmyHCIABuZrXv+YtYAPf905+WpsS2gSQqIhv4V/+MvOLuEKZZ1lpOUi
0kPp4TolVkv6SVgQ90Y5NkCfDj6qEUHxuBaXGM+MSKK1dh1DnYc/dF7L9bos9Vyj+yOgwWKdP9i6
2dunQUZNQ3awwcO5YpIoTnew0Nx+LJ0L368XPg9k/Hm3vr+l+E08WEzRGmyEBXhEOTw1f8VcGg1O
j7Ss01fSNg1cSi02kpF9n1BXeuwr/iouNffZLYa8td6IaT+FjchG4FGZ0x+MZ0dqSKkeRQc/4MwL
Gue05jK+4wgmWlRcdaf7uhHt1++gphA5kdGfgBGuHxxYgjGi8xdVm9JpuJaSWmoLIJgmL2pKf+Cr
RQyMKaEUJSJZrj+cBkXmv6J5VZU0A1ZhY/fB8zG9yDcGrlsLDeBWGQTaxMEtED8PnfjIMLQ7/FpR
RhnFE7ZZfFC1UF+Bv4ed9jeA9ASiyhOeMzIduOCsptpkT2GZqcxDORFj4cHj5X32oKAb/Sy8VzO4
PsUzfbr/assRo/HYSlpNJvYlWwvuk3qCuPWuX1zCwR1ZpYG67ItKxMfaPgw0ClgUdghE9aitMz10
HgBOuqtx1JeccSXd1E278SY158OcD/opFQro7o4j1WknTToqf2/M4qWAWxypIOXCrQXD9g3Nl4Z+
N1AkRvcvEr1tn8kTv1pVJqOX/teiOIC4v7i5AEh0za8e7H/30R4ga998uyw7MwQLrceiYHd6O5oP
25/NcfiRRNffV/JDLDcaRNvkxzUx0v4eBHP7usU51jgPRUT+uB90rxw0VDkGkRsTbOZ9QRiVrmuM
jgf6YjpXkNHcHbBG3csIhFXtBsn62mj9iD43vmvLth4wyEU3/RSVmv7NLgD1trhYE55DcZAXVtfR
iZTW14Q0pdrhBpcfMvD2RcLf/Kxkj0mhlvMtGqg+fLmDdTJ2xzng741Qxkjo+uUdMk8MtD+HezEV
stfr5anCY5sPvZOiRVEDQ17ECCGplUwPjtReCX7g7iCA1SqpNQTdBUA8w9cZIONTYZdL5pRdt/Et
LQjI5AgD9N464nI9/ts/k3MDYdcI5ESaoaKn/IpX3NBrSA6TTFK67D8+Ku+Np33zg3csOtlUnfZa
qY5tHby2ioD7N0Ha//8KNtmJ6vz9Ag1khb2By6/701bRPSLSGKeCKSj9qftQ+RbLXoBX6EC1I34Z
bdFCshkrlxMjpaAkD9KOsWq2Y93xTE0CP6m/V3Ng6CrtMFv7XqM+UPGWBLaS7SJIvpFjsRxNy90R
OLy5FiEMEFkS/SEgr/YgQDatAma74C3IeodvGMpLduwT8tDodSYArCOWVQNUulZtlM0pQHOqJTsV
UsnTNqESgWUd6V1E0QUjiRhGTS9M1Spq+B4jtQrfVmJ/PS1K9Wd64YPGN7zZjWNeNdMVeTL5d8/m
z1V1sdqlInsCy+ClCkXSWe7M6QlpC78YQ0LXLaoMBWj1sssuTQGZbMup+nkuywI5x94xRNLDJNsB
uxIP2kCQuPJNyYGAIQHH2TKKbVzzgkidPcm8Sx/bsRVFpBkb/b2JtcoCmRJgzLmlyxCwFjV4obqO
cmUS/7WkRUZ/6+ncEeUbRY5ZkCHkUD2Zeh5hyqBqcOGGws64+JQuSC7o4ChC0ozor2zKfTe620f/
kfO5VtREqV8EoZpLJtphioJ8UCQKIUWtzOXErIzIbo6v8rBUQ9z3MHTHIqVY0QpA3o8AGJnaB+ip
R3na4TUAZY/Nvu6T8iXEBDrPmUZdxGjb2fHPa8pdoh7htNH4oVkt0J09oDU3sKPP5U2m9OWkRDDr
nVuE/clBRNEsGWZx9J44rC2WZwjs+pWH+H1ntuZ4yrayW7WSnYnxjLVd7tiunYZGA1Hfca2DsaYq
i81yPL1iBE5tmMVrjgYkpLEwVr1rIgvb944oxgaGaWlKm/66yRtDi+RwW4tTzoB7oHG0SKFNooRr
aOU8rpgS1Kxi1BiU5ln01dWcBY4M7eck42q8Rr4K/neZV6M7iR9Llogvu18k6HwxOgC65RvDeiK0
N/iZ/rqdb4D32tdRlTK28sbP4XOHJVD6M40T5Ho5ji4L9O1tXL0Ox0a3B+r4nytEO06LpDtWC3C9
JYQ931FEeG6o0OP30VESOwSMRn3Ul5LLuOGdH1l5oy5RG+P3quRTCEGYLOynkXWrpIXvRGwvZVqF
fVoWfzTrnc7lgI9K9EwXW7qbo4EdnCVk49HS0vJeOHcAOi3HbPdgJZdmNtdUd5exMU0NEi1CXdlN
JGy0cV314Xy277EYt3gA+nYIjc7+AR7hRaVHFVa56DdnX0hoHTZINWBgOC9FZRAley8my/BpxX6d
TyYm3dD0mJQtcSSmG2za2Kmy1PLk0GHIf22kZE3k+o8b4O3z/hF3fgpuRjYxCy2E2misG9Gj6i/H
L7XDRRrLPlZ3wwgymKUe1IQoK8m3lG8vsSpLkhk07VASjY+jVzGajvxSkRuRgxqEpgn7Mfsq4noS
d20MSvRyUA2SAmws9GaqSCs2cRXMlW/EpTF1QbvSt7C5R/uHZCqEJIifx8iy/un52gynSFtnZsjK
flzsMo084qOd3eAb7BnpjhxjU1+z8bI2tMQ6fAc755l2W+4dO4PvBbrBSASgYr7+c4UfaWPMFr4Y
Q98DFv69mesH0V7Myn+u9WbRcFIDsZkYgX2olocq7kLHim1ebzzmXZGZMTYUhlZwEfAO56145ten
GmvsT1su0MlNFdpgLcFLc2UeOF0CV6Hf3LUGiRRxQLAHqxVMXaoyKSSJOoMZtn7sD8hQwVdrqScT
Pvqng3ftMlohXYTxSXBwa7rF/A73aUt657VtHEJa01fq37pvu5T7o7C+61OltYenXpsLhIf5dI6o
gJO0KBcGbbjoO3JeMi4uuQetBhEH5Q9rQCD/dQE2hxeovcp0Ml+ITjdm8M8//Zl4QoPakYyhDHOr
gEpwJLpNuu5BW7jWuwys1PNpnSCu3SXKbjgY8Us1W9r3Riivwphl2eBwkuour+lU8zm6R5kNdDSx
QlLYp5HrS7mNab/1if6p/N+w5ybJKWatlSJ4bSJSWMET3iyiF0ZcvRPUrpdvBa5H3/Rniuc2IkkN
Ra2azULaP+5iW3bLUaR6NkJMWzqW0nmL9B0V4wq2MdndvO5cuJ3OBp8qHUxChl4veEKvB6Fjzji9
+RSBF9287Ez9DlyVTSTZ10W1Fk8tWOM03Ow4I8g1FJGamGBZ4hzxVVUxQCupDGjEqg9tg6dYW5nV
Csu3jXcripxAOIEGyKm8X7Y0hOFMyZpj2CztGQqY00LK1GCsx+iy1vxO8eM/2CFyjPVjpDYsPEMx
u/Kv0wCvWRVg8Z0+0axQeF6g6KzhGAlFPiXUrZsAcA9Cuo794cJxyEE/4iCqQ+DiYGP+NPds+da6
py7iGur8CtQDxN33QFVHFM+/dlCviSz9ppM4UMQjRunmcXP62++blp77dTuHxUSYD6F71YcfrDpJ
pOUWI4QFlmoemqGoPFhNC8DL47UOPHXbWBlsde1vRDa16+5uHbNDGUFraVC0jvbjl0RBtjiNBb4L
foZw55LB3hOCDN6b3j91tUXP0E7uZFEBEzFl3iQc28TJjXSBFWnzP8uZN3tgMClK3rBrUQz3a+th
oYbZMClcv1PGAXppMzOGE7n8w0udtUNlmc4kjID5rEYjS679fEDegxlmg14I2XzCpfkfh1WGDHku
J6QtGcsNqnoiivvIZIZTfjJ/aZ/q9lV+eas5dASZCbse43GXePrD3VAwuin8tt3dr5MPxDOsgWNi
vJGERwpgNCY9KxrJ0QAY7MHi1IBKxIEWsUeOo4Pn+S7FBtFF8yHU5GeQYmKTzKZYmIOgGkUVq12L
yBZG62lGdQ1cMfYmK9yi73/W9yElp2Iga/BJwdwY1+pL1huWvSldT/gZ5MbH7bYF2dV52aINA7jl
bRmPVq3gdOA7tfGZh1avI31w+vpGLyJGEeLA3x2eP8qkcf6rchpzSaMZR8hV1r3r2ZBfTNp2TBI0
bqspTqcez7HNUzB6SnZbKAf5TdCHmiAaCzDoi4CUXtc1Pe7/70TLu1B9DLZwPx5RdYidx/26jQKX
A/8G5wRYKODF8YkTCYNQPk2Y/b0RdGeGd2yez5iut3A6YD0Rv6ko+VBqdkwTJQTqMYHoBR9vASxx
Yiou+rMrVHg3yau+WRwNUDdlt4LlncllVDnKyof1F7KN2A390oRhcuQ/5riFkABp9ol4wDSKaqPl
TiuwTQei4ummqN/AxvRIjSBDYjCdg/xZ5kkWyaV+PSmFv1O2ciF/Dsy9yrGcZnS5LBWXKhe8e2yb
6WTATBTjDceYJQh5TFIzNBQ4rMpWLrjNb6OObUQXgOiBdAoQ/VDZAwyNRLu4zSMay9le8hF4AbT0
23MFtXECJgGeeL8YVoQEPCqzPGp/l9d41I/qUUYkDDfVlXkWrrDDy47Z7Zi4p04KUPav/kHllf0t
eScOUREfSTFkASU2WLqHRRuzIe6CJIxFAHfQnalZB3+byzI9RwUMHdA1bSQQ+toF2ZR1YYMtKnuE
xeUPoSQYA/7rHg8uJpLDEG1q61aBwwmfD3cEvDFRKDne3WqdSwkGTx4ur4JEi5ox0+vAJymyo3FS
6OQpJx2bojSuBqcwIwKthINysat8KxdPX9pVEqjgA2XOxKBA5AyhqS8VCeD0wRViNBvqrr7iltKP
iuWE7UaAQX3LiwkF75TgoTJgsvn4clKDAUrpNzeQK+wTskMVudTHsysQMvjBtTmB9K83oJO+0KVg
JolXL4xphIlDXiSN103GQFemzDxR0YhB4/0xuzBvpgrbb0fC1MGoHd+19EysBGo3fHzsPCPVs05R
rrOnLG72AaPuKjMC3GdgHLFCvQixmpDYy9naojgfYPU2/Qx/f36SGw/7M8b3gt2vHrP4Q8KIVO8n
y5F4X+iBU99B79uFf+2QBEmFAgYvJKr9xvxuvKweRsf4bnktUMZcnECaVd6XJFtwp3HXf2TnYWv7
YPqya7JM1QG/zVPwl1uLnwL5riS5kYe0k7S6KZ6uJ+eMslL1yqRPhoKL50wbTAfm8JEjjeShNOzZ
XZpZHZrLgjzkDv/zOdQX6VFvIo7OwXC89fpq5jn5v8Vg9snSkqA5564MAJ3hhnC0v9/d0RrtOeUb
Z9NPlzq+EQS/YiOaGzfc+zd74BvWJhj9aXLe6EX2hOM2vH5B8hZjCfjJerK5w6s8SbpiyDBB6RAc
9+3rVp18Dr5EyroJWA8S0pw+Q5Fk4KMSxK/ZKDv0YBvyVWDpQMyZfy1BuFJ0Z9DN8xZV3kP/ofcz
j5dW9JzKjn5OxBW3Rsed5jB6lwkcTx5YwaCQrSlNOfuZxIeEXzs42gC6AJNiupZyZFNcyZ+N0XC5
kKITvBiqHBhmEdvKmxtfDsokZ7eEZOlNmu/aJD4H2A7fwFiYnNuLoZhnj7who5PS3UuexnM5Sb+d
lxl/0g1igqUljoUsreCc6aGnr/6RoT3LQl7oGj6S/vXZ7ZKrPLgvkuo6+W9bYQ4BO+i9SEI4OjTY
WCnQ3L6sts2kutUCosCxVxUYD8bokUtbnCOr1mcqpFDb8DwG5p6FVKWlXWuTcqmGpsuWujh4zpZ9
KaNm9vYTH2evqw9UJdz9G8jxWxIV3kB1PNfUODOX3xB++SmPWu8Bfd6O27ToGIHuGmrtPSeQ3l6b
QF1tw6XtJxCWd69u5weVvIkPp0UH/nHz3Vm71ujtgE7Pz2PHOdVvrVE5YS0tqluj6VNAgtAGnUHc
eFMABDue5D0O3NC+u/Y4MgJGctvenHY/FJz2Pcuo+SRqeL97pb4je9ibINqDO/xhcaD+OPl6kd2j
4wtWrzuhvHBkHj42hwe86yEY3hK1Blq6tzgLH9hXMToM5AjHzVXo0mgdvM0PrSfBB2s0Gqd5Eh4+
XWNIkFqGhI2ljPL/WHrsdzMNo71a1wxU8njEv8FineBn7EJeYOzHiSHbqcdqUHxYDTO+ftwqBYZr
dCx5AVnng6tdaj7+1I0Ex9QeBmay/WLakvjyagOEIacU+Poxyj2G9Z5/67SqFWJWfaqA0ZvqKpJI
KO6NQ08fQ9SPUgognuzbyIPmCK/p36j8s/iS9/3p++a1NnA5kHwJL/2SzWDYPAOAs2nKzCkt9lWa
KNf9aas9cGbUvWAZE9DaxdtZVygJZBWcbtopLlMiEp6dYuKOt4v+uOfMGoU/TRWrN4CYoKlh2Zc+
9bK7bLmKRZs6Q/ooJdDmbocmVKVysNV87eT9vG5y0GfcTi8mIq43RlvbW4XC/n5g/6eFGmD4AFeJ
yLs2+AZyiSA9BDAHPbb4hcUHRAOUNRKiS+f3sbINCQQiKGsj/0N2IByfNcEoyLKtAMR4MX5H09xb
/wQ/E/3qmgxYMbc/9I6mlKBT5xb/oqzHDHVaIEYqcNLyHU8kpx7eWcKYuwcizyKr7jTYEfei21VR
e1KsxjeRKzZa8v8hC9XFrMKDd1R8x+qoMGw4eUsmQtUwaAyaE2+n4uIM/c1xRicJ/V/c6KibtLkD
/m2kcGcuvAtpg+JaCPuTRGSyt5L6FzxySHGDDqDOjRDTrTlwrRSrj6+dvzRFIyS4/lCKSi5HNp65
SQaDwm7a2NWaUPW7rU7jPsT7bErPI+r08LXOhJYg0fXczIFE3xGPLOwPlldG/riTILbL8tshmoQv
7ciGL4uTa8BEJ8XrtyOKiJvAJAY6Xns/6SK9lnF2dDHorGw00cIVNUmL2pnwDCk5N8o4PC7xoDU8
cP/CR4jGxRLVO09aaP/YVaBfX9dlx4iQYx00iIOjLTdD3x/7KK4IqPrWTFQLKWSQbRNX5LvIlMDd
pOtttz3mOqFdrzKHMjuhWZ9A2g275eidcXW2lRoVEqRAc4p0TEnaKd3HEnI/9u8wKmQJCvpNo8FQ
sqeefDwIkNBpC07zmK1Nj2ZsBFQT8x6drcdpNRvkq+x8ml+w70xooMoMxrqRsFgft56vGpc5uyMK
k0fBfXhRab/P9ppzmlp/piHTmFPkyj7o5s3Qd4ubaL5Zt1Dwmlx8aaz2OU8NhDb04y4JBs9wME65
quLe3QkqsH79fYgloAl5YeeLIhWQ3LRFj9v5mu44ilzi4OjqflsgtxSetgOC4b7vvq/xBhnu2Yz4
kna+ZIgWML4NrdBhPMyd+68/bEN/I8IGcvhiz1XZforPjwHPWamCR/o/lFK3yvxy03MIjTPGVHNz
aJSK1a4KEVLIce7HrwmxLMvJCGTdiTMLy/hIyGZ7O18d4cH5tODScNdgmcG5eoJrgL0dRO94Esie
CcwbyAY7YzEQw2HJ0c0weGJjaaNS3PWaNY1S29jumbbsOVK+FjGAACaqRXfutsfBrZ56lAsSpcN5
quQG8PqyZtywgcfwXrZEMGK5McOlKz6Bn0QrkA1UQ+1296dSnYdyQayqIz5RnLMxzbW13LIEzT2Z
d5952WGbsNewbIiIGxmjtC/FWWAIEhq5nKcV+SeqrfXzO/luF3fIbqc7EhJ58zwemZ1VlxSAjJeh
dYPuhjqusGeSnzvPlIDBRpyliM6kRAtfnXcxhQImyfiYxEphpMzRdrYNKOwM+10JlTLmFfR+XmVK
lOT/rHx08PfdrKZI3ECYboSrfjVUmSte9GQ+CfnHtTBJW2gKoVSLzAfkcebTcfst7DG1YFm6uejZ
K4OSqR99TYogY8lno2j17T4nhknmVdQ4r5A4GkTCkAbFENtuFMUK3DmOllYdP+Fa5Ds0+Cdtfjeu
tXpsueJbXWY/LZ6uN0sy3i1JW6rl156y4Nuj/ofEjWW0CPPAUn8pBgPzlr9vkmvY5+Vqu8+UeZ3b
8Xk3WS7/6rDvtZttDiBkxm/1LBaaGI8Jw/mZPgRVSHq4ex7Hfug2KsllM8A9tlth3sEhfi37eJp5
AHesM0LK9nmZZE5429a2xUcpbm4SIH5D1MMFLJPoBDPb12kIh8ab/hptQRXx8odImER27/lJLYOg
NixoMdL/0NY5kBtQ9R/wrpOL2iP2PnRnZyERQ/y9YhpNI/9NLqFYRXJH1NaR/DiWxGke7nYljayE
zO/lKhMG3kHzG7N9hdkIX8la8XgRFQtidZHUBvwR3fyfay5ifMg3ekKpP//qMnmhDeAC7SCFfMZ/
cCKemNpmXLvz2ccbgSyQpaOsi1wM9+yyb2R0rRka7/EilerYzN2i0PbHAhMny/LOne+RF+IZiXSV
OgoX4bMfNnrC1oA6UtRvvqlhcg83v2t3vCEkLmm1TJtGurFDxp7IhPvQMxSpNd+2l/OYYGNnMAwE
EapRUBQ/eGm5Z2L2zcsBQIK7VEhc2hoKKRyHWqoXxirkvta8fKc0kAioAOE2Oi5YzXT+dKQ2LisN
/aTiA1FuQWTUOZ9dpQCp4wE2C+jWmXFM0q77683k9bXuQW2Nxd1t2+N9NJcJbcopw955DS5TD8EC
Ha54Yq5gE2tkCGmp8HiyPHIvWIIrACjJLSFs2gquFjIgiKoovkxv8FQ8/hLPl9t/SHHpAzoQt65T
NGLIEG+oGgHjmseCJ1Wor6QU3kSy5y4H8F4mDsIeZcri+INqyvXUYk6nZO8DI/wZgdSgzJi06q9U
4jX2deDwv3ZUUCle8YJKrE8A/QR/NJexZ+Iv8B6L0g8YsM6ADbflFFM7f81F/UkGcHqzchoVsw2f
a41ExkBe9qjBfkCUoDxhXKJ4JXOIT5t6VWy4SVW0C397iZo6QUH3kXkmxb2hAFmLy+ZCvseoTh1A
lSe8F0uKQGPJgscLB8ZhLab8//OAXwIOVZJnToqNTZEajLnA7eotqC5YIflHVgUCjDdR8dBf0dja
0oEPBqIB0UwQn4VBKWaStwE6T6U2cVcPUXu6X/CaipxghC0npDqAb8q869qptJ6QpbhTIGXoaYnG
A6HdPvhNJsmr2ekx3QJUjwN0bnFSrUhingXH/w9q7p+mu8Imy5lErXOC2qETCzO3/b1hsEIB3kdt
9xjXkpI18FQf434/xGArFagtYYd8TN2jsQosDP6/4S9QV9F/oWzngrpmU3KZWveB23cly1X+VUF1
cimRBShryVUshy6wQGWt4JGucXA2KxAadRe/InAaRt21NnKwpfU132NBFjBVEXYLHUtNDrPmKYL1
gxEHt/czlXVGu2H4lQfr7l/5169RGRtsFlblgu8PfX3fW3lamjQEhqSqy/d325rRcSUulHE+lRdG
zLLLrRwuQ+KqArNCrCM9A677eeluLnRe+N5lG0g4NdI4E+obCCWAT2BHmHGiJcdBB1VYd7gLKkcd
SJhq40nQr+PhfvQ9iHjW+2KseFDZXdmAeyaxv3WX+Lzrm/KAr39mYN/0IPtuFrJzg4TUQWd4QFgj
c76iIkMiR2u/vvesmrucUxqdgsIH5vXbfndOvMxIMqDzGhYz3DE7qE3beO+genw5QJDgr+FqBCmF
GaoRs6ouHHA/bAiH/IYaFOvsjT6tATov7DxeGrYJqF5NcoFmLY+6p0lX9m90HUwyE5jNOaBno4dz
PrtrF4XaPUltFLSE7ZFbJVW7frehH0GyBGlThp2H3Vg=
`protect end_protected
