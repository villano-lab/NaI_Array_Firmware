--This example file is for demonstration purpose only. Users must not use this keyfile to encrypt their sources. 
--It is strongly recommonded that users create their own key file to use for encrypting their sources. 
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
t5+vIBVZl21TPq+vETL+74rStkW2VXvhT71/DdFRdGeyN9xPB2fgNz2sFwNeQtqObJBhBAICT1bT
vdL9vIpxXuSIcqpIcTx6eCkGU2LR5NsSnvadgcBWo/W31Zo6y2YSLJv9G9Kvmrnk8kPdxGTIDUL8
D9wn34sa0UuuTa79ILzUDOLHhjbx36brtz7Lv5fSJw6t5MXPBCb0lOvgRmq9jVDdclpnqqKevwq9
DTNfIC9ozyzpCpCtJgiN65N/lVhS/kacAFuUkqrFUAmULgrgs8X2Z9MbMmwuJYVcslmKOqd7BIYX
0cIq3pyWIu/++XB5suh6i5ssEqCpVRgLw0uCsw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="eAlaP92q1ViMpUEO1S4f66NpwxLl4NEvqkafzhs1Pg0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9888)
`protect data_block
Wm9CdS816lI0i/pls6MwMTRwMsd7se/ZEoI3/cdFp+wGzbyOg+BuUCK1TSEO+TZBKuNxyoqIIO+w
FDfNaXrC8TFbnVRPGrvmPx+odyvK+YBlXhJMzl+/s4KO09krEgBK3k2yJxvOnLS6qMFvY/j7Kph5
MZWIRjXbakp8Wcia/3lhquiZaAoDKQbWhOyCjuBXF8C7WEw9EQVw1DTUkKkRuloOWtjgO08x7EJL
ok5TwB/XmsTd03HS9Yg8A39LkX5SbgtmLeogNP/H8fVkrkCUtrv/YQNFgrxqvJUI82cyH1dsUno1
3Gs2FLdD1VS0LayLZawE8okDHYwz9kWawY7rq6UZdhkp3RWiW6LBBy3FOK0gA+uYympc6236z5cz
n81I1qGVLLFbwiu0t2TcI4KUpz8/17oQOjMjnmay6PkABH1psKNIvGpbYy0c2iR8lO228UPGskZL
T095u4GbHCtCBCO4HTZMX4Hs7J8Q9FxgMIPYjQMbNtSOUXc5dB3ctiHMjX+39UXwtvRfl9Rlilg6
ZUtE5B1Vj91YdZjmKQOmuur/HX45gISNqzNyqvCuWiZkCO9sGc5bJdzl6U3MfR4+ZlR4mV6j2pZf
Y6PB3l92fqkNAt6vnz5JO0+Txa7iJJEFPjqZvLqFRlnKDG3TtcsYhb37H9EWpjBKBPFlkoAswlDc
ALeLzydOoLTAUr69DdA/AMerh8Fs9HkkGSG0HGIR8dBOd7565O+m28N1RpOeVUGRYz0jMeniKJZ4
nmhJH7tJScDKs3DMUX6WnDa33yd9E49oD9VE7aANhFT6MDS6mvT5Gtwpt5oMbxKvg7DZg+GEyxvY
npAx6COzaqz0ee/KTSP1pSRk+R0XQDXcH8CXPybtbrk5zS7WKkwM2VUrlg15eDPtJ9ZjuSJR2CV4
gexodPe5HLBLhqfA8jPIq2n5wtiv22yOsCeciziI21ZOpNSX8hrRwVGBaKYAazdi8mp4ZkuKS0ld
Ms0PAeQMqvwi2m252VwcMT3mu9l9FrXHlNdDn4gcbN4RDyiDGkOmOxWHH++vNaK/Raq4s+Gj+Udv
Vycpph2bSv85ZzCqwWYVYdbcdD5jXbDYOdFzyrUvzE24G5efH1yXA+47r2Zs6HTs/aMQ2+hP5gZH
74zul/lJVmOm9GnutgWIXTiUd7WYndllUqJ9RSp8O04nsAPzmM03A3DM3IOog0i2lR6JCUw7WbAW
873eTOzt1GR6LfKzU+UlEyDDR5C1uwPsAG2Ly6rM0SlNtOnC8A51fdOjSKjdR7caUdeteX8oOn//
WBYO0xZfahyovfp1yacYfH47ogOdRaeve0/+2/cW94kDprzbC2qyUp1NUMj9NLrrjqoUvb0TIj6j
wyg3CflEUjT21JlJBvJwo8U01v5DtHzWlu7n2bH+4g+aAImlizahPNjIqVTmmooRCOU0Q6GED8Zj
HYwH7Fnb3jYHBCKszlop+/wwzDcZUCNkzDCS2nlcjJEBHLBLOQerEcuFPqg6lSPuJbRt6dRZtscD
6y/Pznc5ltVF5Y9lUlRGWoa4FDo7t1spiC1r69LIqn1yg136GwFGG1erOdlsk9PnZGkilXKS5CFA
jsUeBgpeoGqTgo43qeVQfx2esQUkvu0KmKCljo7I0OWCztu1SS2DS1w8/6Ku7TawqDj1ssJIneda
ANQBVKow3L90NGL0T5hTh5SqTao8jPdP7JB/O25nNgjr0eUJ06sKa/Wm7Vm9iIALWRyQyeVxjioU
QUBO7d+KhHYfUiSqP1Vm/Z4sVmh6cwOKjWIJbjqeZfnVU2u+Vgdzx7z8MfYQhaBLxYecFelg5n53
9axqSysABJh/xwGm+szdZNAfilLfLkzDptEOVxWKtlSFZ7gw2dGduOG/8hI2EqpT73vgq6tQ6UmF
tlp9qaKqbAHPXuNUncAUEMrLTL/wjq66/qc5SfJqahjE9QEsds1Df2inPe0GIaoG55zx/h5kENGe
jKf+PNoovGgclFNKe3VYplD3FIpwUPRHbw9jTShL06+qrmggJ2/N7QCbt7QL8pU26oMrHG88vH6i
AnpLf+sbPeqWX0USl6OUSzkN8173g5ueI6/OQ+0vNxDZYZyOTrObErSD/f417TIBDuIyt6ZYjWBk
fGrRClKl7zXHN1Wb3fG17xXmfcsjvqigVE2Ev0rnZSypG1K6LXD/+D4doOAAvK9gB3ed9mPlLQSq
lAEXjwfMwmGswSNkqApy76SfwMMQAf83QYFd6JT/x9ncM5DAXnjGFbV5EH+zX4DqLCO3h+DfS7oP
VtRq1nZ+jRKOcsw0sgEcfDSIsBv2qoCbEdQMyinYSAdEoC/qIv9Gacym3ANZ56apgHUmXnl4V78V
5zCcZmKKTSWmJVPe984W1vix4oo+dbAadUXqULYQwifkVupmr5UtFw3TeZf5RCqKQVJpefYo+mTt
rqJwgzfAsGZLbymS2B7zrWJM0/H3Y4LkwDFF0pLlQAx7RiKfxBUETlq4/+tIAsex2ybMPxvmNbpY
XT6pNWM3rFbNxw9aNhYw/fAucd6QPkFGCeDDmJTZMC1XePQLX504xtnzZ1mfyh68MkigBWJhSaMu
ZuLqgSF0M9PoZ9g8j8fYhIn1EvJX/HtpgYx93WusNKg8TaTUgkkwgGorp2fdIpclr4QEJTEt5/SD
L9Z5gT/FGQQtSL/5R4CcdXbvXMc7T/2HpHwoTAUvzf6T7wmgp9/jOPQOFPW2ac12nQvzRrLin53L
5KbzyATPXsm5t9KFD7RddrCcypXjqlZqvMrgJFXsswbYIMUR5qDnSKET7tZD/8gXyS+7oMjqvIwZ
+ZyFATMzuYmk89zC7pRlJHdR13dRaecgIZdBXBdrTLAqlJgumM8VFRCB/ZlX7SVCRSXG3rdaNhmZ
Hk6tE7rblQPkcFrfXE7knshiko0cjC6akFCVO9n6oWip+oaQHjTahXmbRx4CtN2o3VB32zOk20OV
M9O1qroXD89LD+XIe7nXSY4Rq2/SB1Cf2cZZIgQqDY1X5//GenQMGa+P7LMWnBwBrmxbo76NfQxN
KYqSnpOERvuivHmKThSq54dNlMrY2Ur0eOl4RZ7MctzfyQVcyimlCf9RypRZ80xMevWiKHwpzU4+
gElZcgThXD2FdupNy8oRz/rN89Be4mD/EALtDGSV54oBFinaQkfUIk8UUaZazgqfpghMKJHfWxMF
EBgVPdBmLp49fQJdPZl2Mepgy6lUO+JduTPFd+Fh9SpvjEJ8LSMAOg4jnTjx5fjP0sFscRXfW+M4
5jvsNCxudqTbBIr8NkXVS4fwL06CcHScV97d/xF1o5blMp5BYusHrL6LgapytWvhpg2K8ha1RKLn
IAIAu0ZlCg3daodcXMmf6cDDOs921cIvGLS1Ee/TXSm93n2hnq7dVEF7t6q1dP1gEoeYw4ipZe+c
8C+SjQnae7Gsh/umL+hFbMcGvcaEiFh8zNulQrpddkMUGBksbU4CWOZtUJHBhtIyAxNTOCwpQkWQ
RPTi6i6/kpA4IEg7SWLMFR1ao4G1llL8XYZsujVIePZXERZDhNqBzdzaOUDfmnu8ZObfqFGcts7V
+BsRYZDZteONPWUvz8l5xHgUFFLtOFEG7lcoC5PrEzSVmRmTGOw9si7Ov58ijo1IuuS+JuA7aZQm
slTAAwv0fbrbhSJERAdpC1+dCXlBwr+7FGyhBymQx8KehFqf1v9JIYjEYhWyb0epyC2IFSIvQGqR
oR+rXsS8E/Mk+B2FFmEil65CchtFmgHdi2GT20sZIh9Q0kARNT9cEGCgszR9bxZPIbgJwXBOVpyh
BiDNVGyjhE0KdFlKDHF7M7m/PENYFX9oQzr75JS7CfqCS9N0ymY3NMud3eFjcgKyhudOP8JlIKEy
PdqQtS0evg8CxWb+p2fTRBdBnrzVsKSsO9qov2j7OHTIELjeydn811KBqI2ozvGyhPRGIGDjfg7S
hRw76YhXafXkyw4qXUuHLyA4gl8PxqrwksOqtfnYprBNRCwoZdHJuGu+e7OgGOfIYFaElbdwDsy3
heNMr6fugeeszDOx+quRkn3UBMdIguBktWqthvlmnb+uJ3NfC2dzXzpFnfPfNkKyX8bQiIE+X2PK
UpNUgGiLwr+vLJ5LhSHLl26yUeFqWiaMAhPqKAfjOQkxr6rs/V8qD3oDQbPaPzk3dsTdekA6ihCt
rRKTaZ4m0/ShOHsI3mKSCIJ6HY2wFw5oH3NTqxqNSBFOKkxh36FbPnYiu23UT1gPN6XOnfJVBjTd
UcWA/UCVCyXTLyHuhcCTpE2Q5F2CUynNr+6T3emEF/MG2C167e9XsWkNzh+8bogmsftg5Vf/xOBJ
QFsxnWYCtKSH399dgV95msbGlVyZGwAlEnuCZc3nP1VFXYGus0ImaSMLr6gUUcslVrn3MFzCBf5l
k8pI2mX2xklyLL0XgsGkBoVrQQrgZGocbGvJ7Q8aL2/aeAmrR9rxMOEwTtyPxh8HgPSCbkmSyHx8
dgYJVdWsLiN7SouMQqUzQZyCrkfJ7PKoR3ZNJpZys+SZBP+QE+1vn7W5s1iX8/sSlhhe88JKtpWu
GswAQ6naHh19ABsjYTqW6GYoGYd9PU4Z7Tu7U297EbKYrazUYaCxyBj+Zi1RkusW6jmEm/pJrNFf
VbbOWVlqxT+4+9t5RRhAFUzlxAtozp0cYyyJuYKwtXz+b+6eTTv7TJKpZPFe5kRKy3zzg16Gwsq0
UrUZyyajcYOSO2A411kNTLTVBBSoyX7tg3mY2gXMXooAqyiRspbra1U67kcOS5C6sTK39YCUMpDR
n7aBh1wyOzyHsiOK2egobLx07AbklLdazzSxy5CNqXIizDD7+UI8pBiZTZ8GxmJPcl7dj5DpeB5u
C9NdeCPD2QZWanoe3z8zjqTEOOTKLF9Yg15/M5dMNRFM6ys3/t5TeBhnHHsKY8j0aeWDOrT5+Pt5
9hJvE3YgkaaJ9R2zquLQKNjjWNOkCwNWBbMtG746bbGgmdKxXpb6SZP+D8AHSS2ZGyus5V/Pa7vz
DSGpxDDu/UqPRwQDnl9xNc8rxr7R91c328QwhUolCr6tOG/lDVwpIBwlK8ySp9cPFq2xsLj5IvH5
+lKEZHHLCFghQ3ZSKU1dRZVcYx7J6FNxiPH+G2Df5+Y/U5Tb9zX0mHGYYy55ZPgjhtFqjNkO10Po
1/FVKMv2xrAoCsqnVsZFUlkV/M01rbez+zBoLMLvTqtbS+Gdr08gPGuR77BlxsW0NTeHhvY3s4pq
apMoOkJDed6xtTRqoa4c6MABhyI7rH3DmbvdawbGS9ERIP/3xYs1y0W4wGS+AeFm1aIdb4Xg8iR/
bMMWztHsmVMylVu/Im4kGdv6mci5MIjDCYGao3WPFH+VDl9+g+mZxvkRYC+UC9b4K6ZuNaTw600H
pcCl9sVq+Xbddpoturgn/K07tzLFISgVv0BCHzYPH9qpdip2BIgig/gFCSKbFM5V6BHrtm6T0xEO
qu/nyqpe0aVaPlfToCD8dmTjA3x5rus8o/jC80ypsPTF97NRjebaCWqvh7qcKNaAd0yNnFKu+MnW
vv0UFFKJW2QEA2UOdBMy8NpLKgAGK/9N37yPAP1qxS8sSXShu9PMIVM222kRwZDQ+1hYg/nsX36u
wbOWOzzrumFTu2m14+4dg0MVrN9PFu3dWrigNszVe3oJ2jbn5sDgsYW+ZvBBNj+xV+yagjSJzLt5
NDJeRIESdQfXZHjz9Wa9Tw5NAgqmYgHPXy+ShNCsl4dFUoSHzAR4syL4rnq46NKU3WAKJnJeb+Th
HyVWSDwxNP/spHP9lAqhYf/kMiBnJrsr9BPrAiWfjK9tOUZ4BwFEx7FRHD5pmIKVs8ndOTV0KxVr
NAiJ1UDl05rDGUxwM0KGMCGLywWGb2A3mUtjPXq99jYd7WD9oKFTmDJ3Ku6w/kTm2gPHKk7Yv1aB
tIa/bYEyQMDqt0PSc1xyXmWwn//CIUHehwS9+KbQUMB9Pm9/PMegxnTzAoGr2lakexQ2YqcPPLfa
BQqov8a2tqWqQLKPXHve+QegXJC8bdDTlxaK/OuNoyx7t1HAVsPQxr5YRGOz4tw0Qgwh34UXq29p
KFUKOS+77wERoF5LpxV2KSbQS1c37O3g+VVED05O4oQabT6c1NS2dA10XRDHVryn7TL3M6y2MLjR
RjOK4u+15QjMZZnoQU5qpDOokspgxEbub73RshomjEQLbk6SG79VviywnUt5zxTlvPcHPZb66c8z
RwV+eUtcNU8x0oflGmDm6ORpx+pAEaCRtSGmkPg1LCP2ZDJDc3u/NzmAzEa4A3L84i5I9/gH/FcN
As5yo8C/QxUtEDeFjvu+lKIgD3M+7o7mmwgo3riwi+s88TffJ3VJZdnGCb5PGW+CDZp25CMem+zn
CyBU/zjZBlct0idCsexFCfwYJu0hOLa2k5arGk+V2gOlcmcST+Q0Q0cDUTpB5GDC0ONfL7Ka/8el
lUj2pWe5bXyT9C43V0eb5LimSSXKlvTtqc9i+BXAdS2yL2aWmUjjeysq6nS/XRHMVUhXAMGRM104
szSQT2RMNBX8z6IsFBmvSYd2kfrgwx38IByjo88nm4tIf3YjTfYjFaEDql3O4MZYWadcRIN+WlRx
CAFWPZ5LyROu9fcepgvCRFUYh21MFohpg/1BDwQdhKutheqcXziIrUPVG9URBKJ1lZtVKcxeBNmc
DUma1sOubXmE4KTiYq1V4SQgquvWoIPhI/a9JUyElJzhd7hca53lzesrhZhc1WfQlg2OxBQVUcfc
1rjkmWbFN7n6ARlFrzW7fkdG8fYi3xQuMwwKU+dhs9vFKC/mynpxTStW6hHAJUpA4ghgRnk1BArB
Poh6Yb4uzfeF/S4d48EmFuo2yxQkMaJE60Kx4aclDE2bEjbfbOK9oNqKTl107j/jugy6T5K5NR4q
IGpVEVoHsOn0dSyimn4lcOuL8k/6XvvRxbbENL8u7zK4C7v07Bb3QWK94H+3HbupUoflBOOc7USs
P+E0E9gyfrYi9g4+XVsrGJE+Y543MPRBlISip8xoazf5pVTOcgqERFxYomLPIxaXsz8LmPdA5Uix
ssnJIy3KrTDWASNGHEmqRLMLk+sSYxpcX3pUXkQbkDE6d6Ie8WTdpRWuecM7oaqr3xeLIHS7J4Nm
rV/YU5X5cs5RTGSugO9ES/wqlQROORRStkf8oEexTgv5Io1vtxvgNNgerq2bgoMwDv81K9D/x0iV
7C9E+5ffYAHe0ImIIJcV4o/Vp08OZMXcjSd9in7aqzGkJdNs1ta0wWHQ4vsjyHabjljY90T0GEDO
GuiNR/gcd2Y+v1eSZGoJEwlL+pk5dFXULoxe04iMVn6MSr+jOIgI+yjWIAXL90RsQ7IZY8uNvdhb
ZnWUQiiNRXWcqFHFK7HtNLWZNt3/ywyCtdLsxYsq2zPQbIYjnIH4/XK4sNNJe+V7rY4AgnvPAuis
VNxGOprUBOG3M2WD6Ow8n+bByt1vYABNqx+H4EWQ3NFVqx5wM8RVK5iKdXyaEE8B27AYOoF080f8
4ba/dy3tzxRnuPV1Naq8mv8jYZU8H1MMk1yrMcsLwl0JJNTab/p6G5uDe/IJ1c9pbJ+Hf2cpSeYY
TONJa1BinvvF0RsD6rJst78IBRCmwGKENISlqMc57BeafS1tlHOLWqoDwGLS0yAYwzDr0Q/KaJVf
jtv76xgYbmo3Q3i6BdKunjbWlfjWKvMk6qN87GLQkBvsVFwKUMKgP6PdiFlxcVG9XPb009uxPOMr
Yf35/pVosywD4S+UfzxpGTU3y4fRWyLwh+BudWNt5nQ/0T3vvQjIssG3RTSbUhuY5r5QFKsc41DW
Bp6RFMqQydhFKgmRDN+NdzZarqWdZE9zi4eSaV5paFJSi+WCAvkJ45F1qZ3g3UGq4QK2dluwJ74Y
g8CNXL0f/Uolxdc5BCQA6DrmN84DjIoJd2rfc3QkQ2v53erGgRx1c2CPddltMB5MdyFYt4ReoIM0
2Q9gc6oUdpRGLISAjcd9Q4Ro/CpAF+4ZeRFfte941S0lRlPQTbS4d3nYVRY8hNtCXK4xgGqX0Gl/
0NovrECLLa+GnZ2yyEqbxnRY/o0swO5VWAIfqEmy58v2oGOsxoEsG9Srmu0aYFhbXu+B5lKDHmmI
piASsVf1MdiXHdeScqA6LjZr2hu8uC9KAFa0ON5qNTNaJaxJSNFKB/9aeVmtCNyQ76Ll8wt7Be4j
aS+CLUI7G4Mw8M/15xLsNmqX97D3tBBwd+yb3armMWUJmlISg5U4jYbbQo3nsH/2FeoOCYx7DHm6
3y4V1rtsGO74EzZgGGkUmQS64PLQAXgS+COHQTvhWgq+06WXwbSZq0ZJmIruN9ZtvBuDcTD2b35q
c+M2m4EeuqSK4kvxkv6Rd8eOLKIg4toI5dqKcp5NcqaPXAxMYpzc3m8GlWOhkJ098D8Nn3VoIMke
WiuhkuhF9wchvkTrs7BAOWfcFj5KUPwNfhonE0LbZtV1v+sewEko/pMKSTCylNk8kdaIdOGppuJh
TP76F8mlqsszsucJkxSUWeqBEM/67jaaMFPB2hupDKiLZOFdR7QM8yiscxx3gaVzp+neXProOzYk
9xIHh77W1bkcPvslDelwhEixfp1h91eYFf0zZ4Eknep/+SRCc02BmmzmYHgZqrdvmbkFe6v9ofg0
QxUV8jzpedP2qwSX0vhKGrkzO7L6RmSB2VtTXTkYECMMSc7mdxNr7Z2VYct2XKV8/rAs8pXCylj7
61Ud/KXAkGlqPSGc3rdvMCUOnhQbsAnsEY8OfFq2ZTGbacHtGDZkRk8eRsUlwGkY9O0KMNxR0WJc
PKu6Dob13hCgcq/kJhU0UN7fq9L0ii8rHdNsxq/WKr1Gjbat6mm0iXQqyj8neczUTPpwWOMXPRtg
7V3IlIKcALwQ2YV8Y9SHswzfGhgh4Ay+CBlbJkNhWvgj+Zc5fk3S0ak2zyaENndXFh+s6j9oU2fn
nGjwzMhnQ8Jaqxag6+N8ibh/W3vufmqLSbAQf4wVR60LPNBnBIm5ZKPLq9RlEkjaEa5gbJJBaoq2
9FhcvPr3TTNibOqtzah/3h+qkAT7dYWP2LedpDZFfMx5XaaUQZdlcaX8EtSebi3z2GhgPspjBdQF
23i9o3zjWcJ7mDzXvSqS74Do+I/oRs72e22D+FYKWQG76mpvTKRhE8sTJSSIWH9KqoImf08S8sUG
B00OrTNpHQZ50SUUL1E1lnogSxNqocN2Wv0TBsHktsM0wddZf8swiaEdwQR370T0HAr3ssOTJoAN
IgrQm0JqRU9hENa/LDlAn6kNZm5XybN38obsNnlGIWwSY8JNk5QCWfta5yd6pYveitFVw3JwOX4v
VPIJWkwk59JImeA3xlBZd8/vfhcYgUBPIoT9u8e8xUHjOxL6rV8U9L9HGSYtXcgIc3wmUOuG6CG9
FGv6ryB+Y9ZsKVJXefai+KpfttSLBvt5uwiEt1GTZIDZlNwQEFgD0LuPfQzCfQfAYx8pHl/RpIs1
wOcR2QaeGKYbrQoX6DC7i6wxVuVwnO3Ooly30rwRmb0aNOgf7IDLzUtsN93WFji681dbVWituxd5
+kb0BpB+QBx1CyhaE2gWcSYn/BY+uNEE6VFpJeQFtw1XIiDEo9Lxc8yMFiDZ8Bt71DDjkJY1/YDF
uG+BgTL0ZqPu/pZNlxhKusBUR/6wZCctDBC8tBcssokZdXsDL12huKPhjVa9DICdbKC6Zxy5ZVhg
/qOevpWaIk5uRYe7sBuAcMTyczJ53PuMe+EL20CXe70/qHMFSzfEugGRPnDtax0k5zD7ekiZC0OW
IIUSERTj5FxLAe3Ji8G7FfbqLwiEKgrM16NH5pBJR2dMpziclV+eodWxUO1eu8GE/DzNnO7oLoUJ
NN78uF+ij7PKT8NglXzFJN97PCYUHid9zNcxXf3oe9QOLG9ld6zVv11Fs0yL6+eHSJDZ7usRRmD9
ZgFLL5A5ef1Cayvr8JDkF2adD+vXlMeouy71XvftlnISlzQy8PTexBCPfIVMyfljnkgR+f3qe1xv
LRj07+Y4+vVSzWaserpLLK9PPGmjr5pK2PpQTECndVkw/wgRB7naxT76OvIw2XaMGBnb7XImu9E9
P6DHDLIwxBOs8nmkbMgGjZr1SpA90IJxmPpC0jGfWzE3VYay7NykZiwAmvzAPMXYjLWmwJETa2By
SDW1WYipPfvi9tIuWP6ER9yLsJsCL8Q7D6Y7T/IoVgKPO0wg3mYGy7vRWCsU+DKiDUYPjB9fJZ4+
w4Qt9en/CiNrwoTXNbSE3fWwTkXogxjgRVLi81+HX2bOecr0+9GMajaWV1nbqUJ4pXIyz+qOCynp
LwQPN/yN1/EttzKcD4dgusUjZ1VE/FSM5C6SsZK27UEw+YctnD+pILe7yxMOYRWKO+xFgQ36oEby
KNlFUu8zQc1xloPwtoq7cdARpXO0k7h3BdCpJDToISe5GSWdtXpUAURs6fuBMxPfmd6oV8cRmzp8
eIM8vG0cos0lE6gLaNJ7RJmSfunhap7rcrQwCnKtM1gmwbwE/NRInHAHz7aeHKbIwwJxCWVX1dz1
mXBPi86RoRjGrRsao8I8e0EQV94sjD1Ujec1mGYx3d2wlptwvJyZBr7O7WbHzMQ1LBR3HMJmrToR
LU5TGLzYKDyHFd7YlcZVHZQMHNrAz0dQpZXXSaBh3GV1mPL6WgOQ9CLvUeGfi6Nw9g8+6AKrAonv
BDCSJwpHBR7TFbyXFOe3POHy4JYCWRt1EBmgetPrkgrC0ciG1wk5YxZ1J44w6x1xVW84576UNS2s
zfv+dGwKBZMXtzwxxx+dfWxUwiEE0RGAyWNE4hoE9b1hD6T/diMt722F6FAE3XkegRmKF0/JwFNW
cVDrp0lDBC3C6hpeYgGU8VQvmGmc8IADbGRqUm5JJAeSMHnItxx6JjnpdvomahQx9L+i8aHvh1W+
X3bVvjOdw66aV0o8Q4/Z2Cebnyg6DLDR86n5EjQjT+YalbRLTPwjOZCjhtdJQwHmqtgEiJcv0WzF
mXGNO5ZoWoy4L59vKETvSRM1alVLdsggpfq4PayeZkhzl5dyvKILvWOX1WZbWTZ5oGC5WBvQ+g7k
A9mvyxsfu1o+QNSFqcV9t01WKfTF387QLLnHXwWfbc7YK/Dw3uuPWy407LGqSa6Q3YMtkHIAFrog
ZJhtR740bTpfx6UIec2uJKv+Je0d50sfcbPsmegv6eaYfHxBdRaO0QwvnDM5WAKt8mNMIR35qNn8
oLR9szgNgrgd+n+OK1JAQARrbCnAWMPl69IgY1jpT2xc6EiS8MbebwVFRSA4lJ1vBHQqzgEqeNJV
T06c89JnHq5qI5enV4oC0zX35rzpdcDyVtOLKd10PVEysG7lqu+lajch5SnKptG+w6m6dxYHXJqJ
EXA7QE/rOhcUgTBB53Sr1iit5XDVMaDzaq8sAieGOTM+Ub7/kzZfvbnANa6nxEDN0D0i+J7TyqPL
ebHp6OdXlTy1S/OYsnmLX9pLHsrPyZ3j+tEx+zLR9Ou8OTxbitG/kERH4XHGQFpmgh9zgyaou/Y/
qdllTL4y3v0FEUxUVSfRio/wrfU/p9O0wWGGVKXsGrSRDqkaUHQe8GaAejMumtpVebjwUPDwz15T
St0XOMTtdb6jxttIbOarDCnzBQiX1kiJ0Hy0jYhJdvwbqWZy2gSB5Dwvg0sVSi62X2zp9kOzmWSe
7oKzfUl6EEULXNt71KzyHGzFq6GsLRIKBUrKOwO8UEmtiC4XQxoL1cSqniBlZzTMZl5jqvA+Z+1K
wN73WO1Gv+0Qqdo5ewhpkpPiX6naH+JB51n1EJtBaYeEI3NzApZtRY4vogw315xqpPb4bBG64hi9
HbCLbbGSzXvAH5+vSIG6o2OskpfVmZk968skj0pGHudgsRhTbvAohrpEYn+cbid+GLmPYtCSB7T0
W66nOBA4uawoPm3lId76Xaxbyg50WcippbI09aCBjB8l92kJnL8d15CeQyOu9W+OIiK2YOnlEXBs
dmTkqFJtecAUBIJ6v/n5jEDZh27NuiZyYItXqnN7VeLV1u1OhPQ7qoxqRvDT8IJq014djLWgwkmM
UDz5Aj+MSQab6ZsFs+HuSaf2KueVz3hj1jOnUZK0p1jkesPcmuqsqJsai3ouWVmPb2Vc9WqWHtW7
lcZM2leQsGAhaywXlQIkQMYmKkI51lun1rLjC7LrbBLjbgqCOp9YV8P7n451SuhOUO7ryw7LzAiQ
fsQC3toazLHKU+oPGiVZ2OY07mQzZD3V+R/8SiLL/KbXIBX7Dg01Ne4v/SHJ85YBtEQphPO8ad8N
f3ECBBerNzwlYGVzPd6h6f7Yr1Ao6EBRe0NeDVD925pm1ny5rvL3Ai0W8GVN+59DoTGMAbunvjx4
7KlYzXHh1CkwjAKeFLIvKLKUyJaZneed9lX7QZ6Cw5emHyGSfmhT0Ot5v+VKeLjxFX3s5xQfNyA7
9VZZMWcWqiT1cWzZWOapK3GsCfKzNlOXqX+6wcjnvQbTWoALobfHqjkq7n70nEh9Cn99DTT30i6R
pdjhK/SwVrPPqiQfhBfuN/9wZPuNg2cIJ1wHR+9FRYEL1ZofqAA1E+G+J4r531+Wb6wubkb+6mtF
RymCf8lsS65nyD1UVQ4wlhSp8qpruqIqKrxXJ2cR3NQ7C8KDkq3zrErFFc9y4BRq8FD9t4XwI39m
cJxBgkVvpXqvOnGbxcUKTSbd3Oyc8idwOqpuB36HRcqAPoPUtsDLU1M6GgF3HO9IWWXRoL88+OLl
ybZ7vmK3EFy8DRajij9Wodw6dwS0VBMk8Jnx3qHbX1BGQYhapYiauOKBNL8p6yCnUlUoIGjAWbPb
hGqrE3SPInFn5HhcQPc+rk9uLVb6myY9K4owVxjeINBuFC6namitYSjEtlB2ReiIixSZPxuAVQ1m
xXgczSjOcKB5XbAZzAu2oK6oOBcZzVkvb9SNAuAbtFfnnw6bxHkSAqBJOrmSn914l1IB8tQHHs8R
eqoGoK2MsPlU9BwwNtX/yTLNkr6brV3cGGex8aRPT5TIDKYhZdSeOxQVg0x0rL8gYfMonha+WZq5
TAT52Sm9Gb48s2pxnfdZAKI3ObU9zkgdvU2CA8zN/wg88c5HNQmY2brvOiqieyeU9c5HkVEhJM3m
ko2AbcDeYUN85zVW0FFby7jsanwlcedO5ze/
`protect end_protected
